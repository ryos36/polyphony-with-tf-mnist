module do_mnist7_mem
  (
    input wire clk,
(* X_INTERFACE_INFO = "xilinx.com:signal:reset:1.0 rst RST" *)
(* X_INTERFACE_PARAMETER = "POLARITY ACTIVE_HIGH" *)
    input wire rst,
    input wire do_mnist7_mem_ready,
    input wire do_mnist7_mem_accept,
    output reg do_mnist7_mem_valid,
(* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 bram_in CLK" *)
    output wire do_mnist7_in_a_clk,
(* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 bram_in DOUT" *)
    input wire signed [15:0] do_mnist7_mem_in_a_q,
    input wire [10:0] do_mnist7_mem_in_a_len,
(* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 bram_in ADDR" *)
    output wire signed [10:0] do_mnist7_mem_in_a_addr,
(* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 bram_in DIN" *)
    output wire signed [15:0] do_mnist7_mem_in_a_d,
(* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 bram_in WE" *)
    output wire do_mnist7_mem_in_a_we,
(* X_INTERFACE_INFO = "xilinx.com:interface:bram:1.0 bram_in EN" *)
    output wire do_mnist7_mem_in_a_req,

    input wire signed [15:0] do_mnist7_mem_in__mem_q,
    input wire [5:0] do_mnist7_mem_in__mem_len,
    output wire signed [5:0] do_mnist7_mem_in__mem_addr,
    output wire signed [15:0] do_mnist7_mem_in__mem_d,
    output wire do_mnist7_mem_in__mem_we,
    output wire do_mnist7_mem_in__mem_req,
    input wire signed [31:0] do_mnist7_mem_in_lst_len
  );

  //localparams
  localparam do_mnist7_mem_b1_INIT = 0;
  localparam do_mnist7_mem_b1_S0 = 1;
  localparam do_mnist7_mem_b1_S1 = 2;
  localparam do_mnist7_mem_forelse15_FINISH = 3;
  localparam do_mnist7_mem_L1_fortest2_S0 = 4;
  localparam do_mnist7_mem_L1_fortest2_S1 = 5;
  localparam do_mnist7_mem_L1_forbody3_S0 = 6;
  localparam do_mnist7_mem_L1_forbody3_S1 = 7;
  localparam do_mnist7_mem_L1_forbody3_S2 = 8;
  localparam do_mnist7_mem_L1_forbody3_S3 = 9;
  localparam do_mnist7_mem_L1_forelse7_S0 = 10;
  localparam do_mnist7_mem_L1_forelse7_S1 = 11;
  localparam do_mnist7_mem_L2_fortest4_S0 = 12;
  localparam do_mnist7_mem_L2_forbody5_S0 = 13;
  localparam do_mnist7_mem_L2_forbody5_S1 = 14;
  localparam do_mnist7_mem_L2_ifthen24_S0 = 15;
  localparam do_mnist7_mem_L2_ifelse27_S0 = 16;
  localparam do_mnist7_mem_L2_ifthen28_S0 = 17;
  localparam do_mnist7_mem_L2_ifelse29_S0 = 18;
  localparam do_mnist7_mem_L2_ifthen32_S0 = 19;
  localparam do_mnist7_mem_L2_ifelse33_S0 = 20;
  localparam do_mnist7_mem_L2_ifthen34_S0 = 21;
  localparam do_mnist7_mem_L2_ifelse49_S0 = 22;
  localparam do_mnist7_mem_L2_ifthen36_S0 = 23;
  localparam do_mnist7_mem_L2_b114_S0 = 24;
  localparam do_mnist7_mem_L2_ifthen50_S0 = 25;
  localparam do_mnist7_mem_L2_ifelse51_S0 = 26;
  localparam do_mnist7_mem_L2_b43_S0 = 27;
  localparam do_mnist7_mem_L2_b43_S1 = 28;
  localparam do_mnist7_mem_L2_ifthen53_S0 = 29;
  localparam do_mnist7_mem_L2_b115_S0 = 30;
  localparam do_mnist7_mem_L2_b59_S0 = 31;
  localparam do_mnist7_mem_L2_b59_S1 = 32;
  localparam do_mnist7_mem_L2_ifthen46_S0 = 33;
  localparam do_mnist7_mem_L2_exit39_S0 = 34;
  localparam do_mnist7_mem_L2_ifthen62_S0 = 35;
  localparam do_mnist7_mem_L2_exit56_S0 = 36;
  localparam do_mnist7_mem_L2_b41_S0 = 37;
  localparam do_mnist7_mem_L2_exit25_S0 = 38;
  localparam do_mnist7_mem_L2_exit25_S1 = 39;
  localparam do_mnist7_mem_L3_fortest60_S0 = 40;
  localparam do_mnist7_mem_L3_forbody61_S0 = 41;
  localparam do_mnist7_mem_L3_ifelse63_S0 = 42;
  localparam do_mnist7_mem_L3_ifelse63_S1 = 43;
  localparam do_mnist7_mem_L4_fortest44_S0 = 44;
  localparam do_mnist7_mem_L4_forbody45_S0 = 45;
  localparam do_mnist7_mem_L4_ifelse47_S0 = 46;
  localparam do_mnist7_mem_L4_ifelse47_S1 = 47;
  localparam do_mnist7_mem_L5_fortest12_S0 = 48;
  localparam do_mnist7_mem_L5_forbody13_S0 = 49;
  localparam do_mnist7_mem_L5_forbody13_S1 = 50;
  localparam do_mnist7_mem_L5_ifthen73_S0 = 51;
  localparam do_mnist7_mem_L5_ifelse75_S0 = 52;
  localparam do_mnist7_mem_L5_ifthen76_S0 = 53;
  localparam do_mnist7_mem_L5_ifelse77_S0 = 54;
  localparam do_mnist7_mem_L5_ifthen80_S0 = 55;
  localparam do_mnist7_mem_L5_ifelse81_S0 = 56;
  localparam do_mnist7_mem_L5_ifthen82_S0 = 57;
  localparam do_mnist7_mem_L5_ifelse97_S0 = 58;
  localparam do_mnist7_mem_L5_ifthen84_S0 = 59;
  localparam do_mnist7_mem_L5_b117_S0 = 60;
  localparam do_mnist7_mem_L5_ifthen98_S0 = 61;
  localparam do_mnist7_mem_L5_ifelse99_S0 = 62;
  localparam do_mnist7_mem_L5_b91_S0 = 63;
  localparam do_mnist7_mem_L5_b91_S1 = 64;
  localparam do_mnist7_mem_L5_ifthen101_S0 = 65;
  localparam do_mnist7_mem_L5_b118_S0 = 66;
  localparam do_mnist7_mem_L5_b107_S0 = 67;
  localparam do_mnist7_mem_L5_b107_S1 = 68;
  localparam do_mnist7_mem_L5_ifthen94_S0 = 69;
  localparam do_mnist7_mem_L5_exit87_S0 = 70;
  localparam do_mnist7_mem_L5_ifthen110_S0 = 71;
  localparam do_mnist7_mem_L5_exit104_S0 = 72;
  localparam do_mnist7_mem_L5_b89_S0 = 73;
  localparam do_mnist7_mem_L5_exit74_S0 = 74;
  localparam do_mnist7_mem_L5_exit74_S1 = 75;
  localparam do_mnist7_mem_L6_fortest108_S0 = 76;
  localparam do_mnist7_mem_L6_forbody109_S0 = 77;
  localparam do_mnist7_mem_L6_ifelse111_S0 = 78;
  localparam do_mnist7_mem_L6_ifelse111_S1 = 79;
  localparam do_mnist7_mem_L7_fortest92_S0 = 80;
  localparam do_mnist7_mem_L7_forbody93_S0 = 81;
  localparam do_mnist7_mem_L7_ifelse95_S0 = 82;
  localparam do_mnist7_mem_L7_ifelse95_S1 = 83;

  localparam do_mnist7_mem_L2_forbody5_S1_MUL = 84;
  
  //signals: 
  wire        [15:0] add_result26;
  wire        [15:0] add_result27;
  wire        [15:0] add_result2_inl17;
  wire        [15:0] add_result2_inl18;
  reg        [31:0] array630 [0:9];
  wire        [15:0] b_e_inl22;
  wire        [15:0] b_e_inl24;
  wire        [15:0] b_e_inl2_inl13;
  wire        [15:0] b_e_inl2_inl15;
  wire        [7:0] b_inl1_inl24;
  wire        [7:0] b_inl1_inl2_inl15;
  wire        [15:0] b_inl24;
  wire        [15:0] b_inl2_inl15;
  wire        [7:0] b_inl2_inl24;
  wire        [7:0] b_inl2_inl2_inl15;
  wire        [15:0] b_n_inl2;
  wire        [15:0] b_n_inl2_inl1;
  wire b_sign_inl24;
  wire b_sign_inl2_inl15;
  wire c1195;
  wire c1196;
  wire c1197;
  wire c1198;
  wire c1199;
  wire c1200;
  wire c1201;
  wire c1202;
  wire c1203;
  wire c1204;
  wire c1205;
  wire c1206;
  wire c1207;
  wire c1208;
  wire c1209;
  wire c1210;
  wire c1211;
  wire c1212;
  wire c1213;
  wire c1214;
  wire c1215;
  wire c1216;
  wire c1217;
  wire c1218;
  wire c1219;
  wire c1220;
  wire c1221;
  wire c1222;
  wire c1223;
  wire c1224;
  wire c1225;
  wire c1226;
  wire c1227;
  wire c1228;
  wire c1229;
  wire c1230;
  wire c1231;
  wire c1232;
  wire c1233;
  wire c1234;
  wire c1235;
  wire c1236;
  wire c1237;
  wire c1238;
  wire c1239;
  wire c1240;
  wire c1241;
  wire c1242;
  wire c1243;
  wire c1244;
  wire c1245;
  wire c1246;
  wire c1247;
  wire c1248;
  wire c1249;
  wire c1250;
  wire c1251;
  wire c1252;
  wire c1253;
  wire c1254;
  wire c1255;
  wire c1256;
  wire c1257;
  wire c1258;
  wire c1259;
  wire c1260;
  wire c1261;
  wire c1262;
  wire c1263;
  wire c1264;
  wire c1265;
  wire c1266;
  wire c1267;
  wire c1268;
  wire c1269;
  wire c1677;
  wire c1678;
  wire c1679;
  wire c1680;
  wire c1681;
  wire c1682;
  wire c1683;
  wire c1684;
  wire c1685;
  wire c1686;
  wire c1687;
  wire c1688;
  wire c1689;
  wire c1690;
  wire c1691;
  wire c1692;
  wire c1693;
  wire c1694;
  wire c1695;
  wire c1696;
  wire c1697;
  wire c1698;
  wire c1699;
  wire c1700;
  wire c1701;
  wire c1702;
  wire c1703;
  wire c1704;
  wire c1705;
  wire c1706;
  wire c1707;
  wire c1708;
  wire c1709;
  wire c1710;
  wire c1711;
  wire c1712;
  wire c1713;
  wire c1714;
  wire c1715;
  wire c1716;
  wire c1717;
  wire c1718;
  wire c1719;
  wire c1720;
  wire c1721;
  wire c1722;
  wire c1723;
  wire c1724;
  wire c1725;
  wire c558_inl2;
  wire c558_inl2_inl1;
  wire c559_inl2;
  wire c559_inl2_inl1;
  wire c566_inl2;
  wire c566_inl2_inl1;
  wire c567_inl2;
  wire c567_inl2_inl1;
  wire c568_inl2;
  wire c568_inl2_inl1;
  wire c576_inl2;
  wire c576_inl2_inl1;
  wire c581_inl1_inl2;
  wire c581_inl1_inl2_inl1;
  wire c581_inl2_inl2;
  wire c581_inl2_inl2_inl1;
  wire c582_inl1_inl2;
  wire c582_inl1_inl2_inl1;
  wire c582_inl2_inl2;
  wire c582_inl2_inl2_inl1;
  wire c583_inl1_inl2;
  wire c583_inl1_inl2_inl1;
  wire c583_inl2_inl2;
  wire c583_inl2_inl2_inl1;
  wire c584_inl1_inl2;
  wire c584_inl1_inl2_inl1;
  wire c584_inl2_inl2;
  wire c584_inl2_inl2_inl1;
  wire c585_inl1_inl2;
  wire c585_inl1_inl2_inl1;
  wire c585_inl2_inl2;
  wire c585_inl2_inl2_inl1;
  wire c586_inl1_inl2;
  wire c586_inl1_inl2_inl1;
  wire c586_inl2_inl2;
  wire c586_inl2_inl2_inl1;
  wire c587_inl1_inl2;
  wire c587_inl1_inl2_inl1;
  wire c587_inl2_inl2;
  wire c587_inl2_inl2_inl1;
  wire c588_inl1_inl2;
  wire c588_inl1_inl2_inl1;
  wire c588_inl2_inl2;
  wire c588_inl2_inl2_inl1;
  wire c591_inl1_inl2;
  wire c591_inl1_inl2_inl1;
  wire c591_inl2_inl2;
  wire c591_inl2_inl2_inl1;
  wire c597_inl1_inl2;
  wire c597_inl1_inl2_inl1;
  wire c597_inl2_inl2;
  wire c597_inl2_inl2_inl1;
  wire c599_inl1_inl2;
  wire c599_inl1_inl2_inl1;
  wire c599_inl2_inl2;
  wire c599_inl2_inl2_inl1;
  wire c605;
  wire c606;
  wire c611;
  wire c615_inl1_inl1;
  wire c616_inl1_inl1;
  wire c625_inl1_inl1;
  wire c643_inl1_inl2;
  wire c643_inl1_inl2_inl1;
  wire c643_inl2_inl2;
  wire c643_inl2_inl2_inl1;
  wire c644_inl1_inl2;
  wire c644_inl1_inl2_inl1;
  wire c644_inl2_inl2;
  wire c644_inl2_inl2_inl1;
  wire        [15:0] d_inl2;
  wire        [15:0] d_inl2_inl1;
  wire        [7:0] e_inl1_inl13;
  wire        [7:0] e_inl1_inl14;
  wire        [7:0] e_inl1_inl15;
  wire        [7:0] e_inl1_inl2;
  wire        [7:0] e_inl1_inl2_inl1;
  wire        [7:0] e_inl2_inl2;
  wire        [7:0] e_inl2_inl2_inl1;
  wire        [15:0] mul_result1_inl16;
  wire        [7:0] new_b_n_inl2;
  wire        [7:0] new_b_n_inl2_inl1;
  reg        [15:0] new_n_inl1_inl13;
  wire        [15:0] new_n_inl1_inl14;
  wire        [15:0] new_n_inl1_inl15;
  wire        [15:0] new_n_inl1_inl16;
  wire        [15:0] new_n_inl1_inl17;
  wire        [8:0] rv_n_inl1_inl22;
  wire        [8:0] rv_n_inl1_inl23;
  wire        [8:0] rv_n_inl1_inl24;
  wire        [8:0] rv_n_inl1_inl25;
  wire        [8:0] rv_n_inl1_inl27;
  wire        [8:0] rv_n_inl1_inl2_inl13;
  wire        [8:0] rv_n_inl1_inl2_inl14;
  wire        [8:0] rv_n_inl1_inl2_inl15;
  wire        [8:0] rv_n_inl1_inl2_inl16;
  wire        [8:0] rv_n_inl1_inl2_inl18;
  wire        [8:0] rv_n_inl2_inl22;
  wire        [8:0] rv_n_inl2_inl23;
  wire        [8:0] rv_n_inl2_inl24;
  wire        [8:0] rv_n_inl2_inl25;
  wire        [8:0] rv_n_inl2_inl27;
  wire        [8:0] rv_n_inl2_inl2_inl13;
  wire        [8:0] rv_n_inl2_inl2_inl14;
  wire        [8:0] rv_n_inl2_inl2_inl15;
  wire        [8:0] rv_n_inl2_inl2_inl16;
  wire        [8:0] rv_n_inl2_inl2_inl18;
  wire        [15:0] s_inl1_inl1;
  wire        [31:0] t560_inl2;
  wire        [31:0] t560_inl2_inl1;
  wire        [31:0] t562_inl2;
  wire        [31:0] t562_inl2_inl1;
  wire        [31:0] t564_inl2;
  wire        [15:0] t564_inl2_inl1;
  wire        [31:0] t565_inl2;
  wire        [31:0] t565_inl2_inl1;
  wire        [15:0] t569_inl2;
  wire        [15:0] t569_inl2_inl1;
  wire        [15:0] t570_inl2;
  wire        [15:0] t570_inl2_inl1;
  wire        [15:0] t573_inl2;
  wire        [15:0] t573_inl2_inl1;
  wire        [15:0] t574_inl2;
  wire        [15:0] t574_inl2_inl1;
  wire        [31:0] t575_inl2;
  wire        [31:0] t575_inl2_inl1;
  wire        [15:0] t577_inl2;
  wire        [15:0] t577_inl2_inl1;
  wire        [31:0] t589_inl1_inl2;
  wire        [31:0] t589_inl1_inl2_inl1;
  wire        [31:0] t589_inl2_inl2;
  wire        [31:0] t589_inl2_inl2_inl1;
  wire        [31:0] t593_inl1_inl2;
  wire        [31:0] t593_inl1_inl2_inl1;
  wire        [31:0] t593_inl2_inl2;
  wire        [31:0] t593_inl2_inl2_inl1;
  wire        [31:0] t594_inl1_inl2;
  wire        [31:0] t594_inl1_inl2_inl1;
  wire        [31:0] t594_inl2_inl2;
  wire        [31:0] t594_inl2_inl2_inl1;
  wire        [31:0] t596_inl1_inl2;
  wire        [31:0] t596_inl1_inl2_inl1;
  wire        [31:0] t596_inl2_inl2;
  wire        [31:0] t596_inl2_inl2_inl1;
  wire        [8:0] t598_inl1_inl2;
  wire        [8:0] t598_inl1_inl2_inl1;
  wire        [8:0] t598_inl2_inl2;
  wire        [8:0] t598_inl2_inl2_inl1;
  wire        [31:0] t601_inl1_inl2;
  wire        [31:0] t601_inl1_inl2_inl1;
  wire        [31:0] t601_inl2_inl2;
  wire        [31:0] t601_inl2_inl2_inl1;
  wire        [31:0] t602_inl1_inl2;
  wire        [31:0] t602_inl1_inl2_inl1;
  wire        [31:0] t602_inl2_inl2;
  wire        [31:0] t602_inl2_inl2_inl1;
  wire        [31:0] t604_inl1_inl2;
  wire        [31:0] t604_inl1_inl2_inl1;
  wire        [31:0] t604_inl2_inl2;
  wire        [31:0] t604_inl2_inl2_inl1;
  wire        [31:0] t608;
  wire        [31:0] t613;
  wire        [15:0] t617_inl1_inl1;
  wire        [31:0] t618_inl1_inl1;
  wire        [15:0] t619_inl1_inl1;
  wire        [15:0] t620_inl1_inl1;
  wire        [15:0] t621_inl1_inl1;
  wire        [15:0] t622_inl1_inl1;
  wire        [15:0] t623_inl1_inl1;
  wire        [15:0] t624_inl1_inl1;
  wire        [31:0] t626_inl1_inl1;
  wire        [31:0] t627_inl1_inl1;
  wire        [15:0] t628_inl1_inl1;
  wire        [15:0] t629_inl1_inl1;
  wire        [15:0] w_e_inl1_inl1;
  wire        [15:0] w_n_inl1_inl1;
  wire        [15:0] x_e_inl1_inl1;
  wire        [15:0] x_e_inl22;
  wire        [15:0] x_e_inl24;
  wire        [15:0] x_e_inl2_inl13;
  wire        [15:0] x_e_inl2_inl15;
  wire        [7:0] x_inl1_inl24;
  wire        [7:0] x_inl1_inl2_inl15;
  wire        [15:0] x_inl24;
  wire        [15:0] x_inl2_inl15;
  wire        [7:0] x_inl2_inl24;
  wire        [7:0] x_inl2_inl2_inl15;
  wire        [15:0] x_n_inl1_inl1;
  wire        [15:0] x_n_inl2;
  wire        [15:0] x_n_inl2_inl1;
  wire x_sign_inl1_inl24;
  wire x_sign_inl1_inl2_inl15;
  wire x_sign_inl24;
  wire x_sign_inl2_inl15;
  wire x_sign_inl2_inl24;
  wire x_sign_inl2_inl2_inl15;
  wire        [15:0] x_w_inl1_inl1;
  reg        [6:0] do_mnist7_mem_state;
  reg        [8:0] rv_n_inl1_inl26;
  reg        [8:0] rv_n_inl1_inl2_inl17;
  reg        [8:0] rv_n_inl2_inl26;
  reg        [8:0] rv_n_inl2_inl2_inl17;
  reg        [31:0] t609;
  reg        [31:0] t612;
  reg        [15:0] x;
  wire signed [31:0] i3;
  wire signed [31:0] i_inl1_inl24;
  wire signed [31:0] i_inl1_inl2_inl15;
  wire signed [31:0] i_inl2_inl24;
  wire signed [31:0] i_inl2_inl2_inl15;
  wire signed [31:0] j4;
  wire signed [31:0] j7;
  wire signed [31:0] rv_inl24;
  wire signed [31:0] rv_inl2_inl15;
  wire signed [31:0] sub_add_result1_inl22;
  wire signed [31:0] sub_add_result1_inl23;
  wire signed [31:0] sub_add_result1_inl25;
  wire signed [31:0] sub_add_result1_inl2_inl13;
  wire signed [31:0] sub_add_result1_inl2_inl14;
  wire signed [31:0] sub_add_result1_inl2_inl16;
  wire signed [31:0] sub_add_result2_inl22;
  wire signed [31:0] sub_add_result2_inl23;
  wire signed [31:0] sub_add_result2_inl25;
  wire signed [31:0] sub_add_result2_inl2_inl13;
  wire signed [31:0] sub_add_result2_inl2_inl14;
  wire signed [31:0] sub_add_result2_inl2_inl16;
  wire signed [31:0] t561_inl2;
  wire signed [31:0] t561_inl2_inl1;
  wire signed [31:0] t563_inl2;
  wire signed [31:0] t563_inl2_inl1;
  wire signed [31:0] t571_inl2;
  wire signed [31:0] t571_inl2_inl1;
  wire signed [31:0] t572_inl2;
  wire signed [31:0] t572_inl2_inl1;
  wire signed [31:0] t590_inl1_inl2;
  wire signed [31:0] t590_inl1_inl2_inl1;
  wire signed [31:0] t590_inl2_inl2;
  wire signed [31:0] t590_inl2_inl2_inl1;
  wire signed [31:0] t592_inl1_inl2;
  wire signed [31:0] t592_inl1_inl2_inl1;
  wire signed [31:0] t592_inl2_inl2;
  wire signed [31:0] t592_inl2_inl2_inl1;
  wire signed [31:0] t595_inl1_inl2;
  wire signed [31:0] t595_inl1_inl2_inl1;
  wire signed [31:0] t595_inl2_inl2;
  wire signed [31:0] t595_inl2_inl2_inl1;
  wire signed [31:0] t600_inl1_inl2;
  wire signed [31:0] t600_inl1_inl2_inl1;
  wire signed [31:0] t600_inl2_inl2;
  wire signed [31:0] t600_inl2_inl2_inl1;
  wire signed [31:0] t603_inl1_inl2;
  wire signed [31:0] t603_inl1_inl2_inl1;
  wire signed [31:0] t603_inl2_inl2;
  wire signed [31:0] t603_inl2_inl2_inl1;
  wire signed [31:0] t607;
  wire signed [31:0] xi3;
  reg signed [31:0] i2;
  reg signed [31:0] i_inl1_inl23;
  reg signed [31:0] i_inl1_inl2_inl14;
  reg signed [31:0] i_inl2_inl23;
  reg signed [31:0] i_inl2_inl2_inl14;
  reg signed [31:0] j3;
  reg signed [31:0] j6;
  reg signed [31:0] lst_len;
  reg signed [31:0] xi2;
  //signals: _mem
  wire        [5:0] _mem_len;
  wire        [15:0] _mem_q;
  reg        [5:0] _mem_addr;
  reg        [15:0] _mem_d;
  reg _mem_req;
  reg _mem_we;
  //signals: a
  wire        [10:0] a_len;
  wire        [15:0] a_q;
  reg        [10:0] a_addr;
  reg        [15:0] a_d;
  reg a_req;
  reg a_we;
  //combinations: 

  assign do_mnist7_in_a_clk = clk;

  assign add_result26 = rv_inl24;
  assign add_result27 = c1198 ? t613 : c1202 ? t612 : c1208 ? x_inl24 : c1218 ? x_inl24 : (c1255 || c1256) ? add_result26 : 'bz;
  assign add_result2_inl17 = rv_inl2_inl15;
  assign add_result2_inl18 = c1210 ? t609 : c1214 ? mul_result1_inl16 : c1229 ? x_inl2_inl15 : c1240 ? x_inl2_inl15 : (c1268 || c1269) ? add_result2_inl17 : 'bz;
  assign b_e_inl22 = (t565_inl2 & 255);
  assign b_e_inl24 = c1206 ? x_e_inl22 : (c1203 && !c566_inl2) ? b_e_inl22 : 'bz;
  assign b_e_inl2_inl13 = (t565_inl2_inl1 & 255);
  assign b_e_inl2_inl15 = c1220 ? x_e_inl2_inl13 : (c1215 && !c566_inl2_inl1) ? b_e_inl2_inl13 : 'bz;
  assign b_inl1_inl24 = c1217 ? t569_inl2 : (c1212 && c644_inl1_inl2) ? t570_inl2 : 'bz;
  assign b_inl1_inl2_inl15 = c1239 ? t569_inl2_inl1 : (c1233 && c644_inl1_inl2_inl1) ? t570_inl2_inl1 : 'bz;
  assign b_inl24 = c1206 ? t612 : (c1203 && !c566_inl2) ? t613 : 'bz;
  assign b_inl2_inl15 = c1220 ? mul_result1_inl16 : (c1215 && !c566_inl2_inl1) ? t609 : 'bz;
  assign b_inl2_inl24 = c1224 ? t577_inl2 : (c1219 && c644_inl2_inl2) ? new_b_n_inl2 : 'bz;
  assign b_inl2_inl2_inl15 = c1249 ? t577_inl2_inl1 : (c1241 && c644_inl2_inl2_inl1) ? new_b_n_inl2_inl1 : 'bz;
  assign b_n_inl2 = (b_inl24 & 127);
  assign b_n_inl2_inl1 = (b_inl2_inl15 & 127);
  assign b_sign_inl24 = c1206 ? t561_inl2 : (c1203 && !c566_inl2) ? t563_inl2 : 'bz;
  assign b_sign_inl2_inl15 = c1220 ? t561_inl2_inl1 : (c1215 && !c566_inl2_inl1) ? t563_inl2_inl1 : 'bz;
  assign c1195 = (c605 && c606);
  assign c1196 = (c1195 && c615_inl1_inl1);
  assign c1197 = (c1195 && !c615_inl1_inl1);
  assign c1198 = (c611 && c558_inl2);
  assign c1199 = (c611 && !c558_inl2);
  assign c1200 = (c1197 && c616_inl1_inl1);
  assign c1201 = (c1197 && !c616_inl1_inl1);
  assign c1202 = (c1199 && c559_inl2);
  assign c1203 = (c1199 && !c559_inl2);
  assign c1204 = (c1201 && c625_inl1_inl1);
  assign c1205 = (c1201 && !c625_inl1_inl1);
  assign c1206 = (c1203 && c566_inl2);
  assign c1207 = (c1203 && !c566_inl2);
  assign c1208 = ((c1207 || c1206) && c567_inl2);
  assign c1209 = ((c1207 || c1206) && !c567_inl2);
  assign c1210 = (c1195 && c558_inl2_inl1);
  assign c1211 = (c1195 && !c558_inl2_inl1);
  assign c1212 = (c1209 && c568_inl2);
  assign c1213 = (c1209 && !c568_inl2);
  assign c1214 = (c1211 && c559_inl2_inl1);
  assign c1215 = (c1211 && !c559_inl2_inl1);
  assign c1216 = (c1212 && c587_inl1_inl2);
  assign c1217 = (c1212 && c643_inl1_inl2);
  assign c1218 = (c1213 && c576_inl2);
  assign c1219 = (c1213 && !c576_inl2);
  assign c1220 = (c1215 && c566_inl2_inl1);
  assign c1221 = (c1216 && c591_inl1_inl2);
  assign c1222 = (c1212 && c644_inl1_inl2);
  assign c1223 = (c1219 && c587_inl2_inl2);
  assign c1224 = (c1219 && c643_inl2_inl2);
  assign c1225 = (c1215 && !c566_inl2_inl1);
  assign c1226 = (c1216 && !c591_inl1_inl2);
  assign c1227 = (c1223 && c591_inl2_inl2);
  assign c1228 = (c1219 && c644_inl2_inl2);
  assign c1229 = ((c1225 || c1220) && c567_inl2_inl1);
  assign c1230 = ((c1225 || c1220) && !c567_inl2_inl1);
  assign c1231 = ((c1222 || c1217) && c597_inl1_inl2);
  assign c1232 = (c1223 && !c591_inl2_inl2);
  assign c1233 = (c1230 && c568_inl2_inl1);
  assign c1234 = (c1230 && !c568_inl2_inl1);
  assign c1235 = (c1231 && c599_inl1_inl2);
  assign c1236 = (c1231 && !c599_inl1_inl2);
  assign c1237 = ((c1228 || c1224) && c597_inl2_inl2);
  assign c1238 = (c1233 && c587_inl1_inl2_inl1);
  assign c1239 = (c1233 && c643_inl1_inl2_inl1);
  assign c1240 = (c1234 && c576_inl2_inl1);
  assign c1241 = (c1234 && !c576_inl2_inl1);
  assign c1242 = (c1226 || c1221);
  assign c1243 = (c1222 || c1217);
  assign c1244 = (c1237 && c599_inl2_inl2);
  assign c1245 = (c1237 && !c599_inl2_inl2);
  assign c1246 = (c1238 && c591_inl1_inl2_inl1);
  assign c1247 = (c1233 && c644_inl1_inl2_inl1);
  assign c1248 = (c1241 && c587_inl2_inl2_inl1);
  assign c1249 = (c1241 && c643_inl2_inl2_inl1);
  assign c1250 = (c1232 || c1227);
  assign c1251 = (c1228 || c1224);
  assign c1252 = (c1238 && !c591_inl1_inl2_inl1);
  assign c1253 = (c1248 && c591_inl2_inl2_inl1);
  assign c1254 = (c1241 && c644_inl2_inl2_inl1);
  assign c1255 = ((c1242 || c1243) || c1235);
  assign c1256 = ((c1250 || c1251) || c1244);
  assign c1257 = ((c1247 || c1239) && c597_inl1_inl2_inl1);
  assign c1258 = (c1248 && !c591_inl2_inl2_inl1);
  assign c1259 = (c1257 && c599_inl1_inl2_inl1);
  assign c1260 = (c1257 && !c599_inl1_inl2_inl1);
  assign c1261 = ((c1254 || c1249) && c597_inl2_inl2_inl1);
  assign c1262 = (c1252 || c1246);
  assign c1263 = (c1247 || c1239);
  assign c1264 = (c1261 && c599_inl2_inl2_inl1);
  assign c1265 = (c1261 && !c599_inl2_inl2_inl1);
  assign c1266 = (c1258 || c1253);
  assign c1267 = (c1254 || c1249);
  assign c1268 = ((c1262 || c1263) || c1259);
  assign c1269 = ((c1266 || c1267) || c1264);
  assign c1677 = (c605 && c606);
  assign c1678 = (c611 && c558_inl2);
  assign c1679 = (c611 && !c558_inl2);
  assign c1680 = (c1677 && c558_inl2_inl1);
  assign c1681 = (c1677 && !c558_inl2_inl1);
  assign c1682 = (c1679 && c559_inl2);
  assign c1683 = (c1679 && !c559_inl2);
  assign c1684 = (c1681 && c559_inl2_inl1);
  assign c1685 = (c1681 && !c559_inl2_inl1);
  assign c1686 = (c1683 && c567_inl2);
  assign c1687 = (c1683 && !c567_inl2);
  assign c1688 = (c1685 && c567_inl2_inl1);
  assign c1689 = (c1685 && !c567_inl2_inl1);
  assign c1690 = (c1687 && c568_inl2);
  assign c1691 = (c1687 && !c568_inl2);
  assign c1692 = (c1689 && c568_inl2_inl1);
  assign c1693 = (c1689 && !c568_inl2_inl1);
  assign c1694 = (c1690 && c587_inl1_inl2);
  assign c1695 = (c1690 && !c587_inl1_inl2);
  assign c1696 = (c1691 && c576_inl2);
  assign c1697 = (c1691 && !c576_inl2);
  assign c1698 = (c1692 && c587_inl1_inl2_inl1);
  assign c1699 = (c1692 && !c587_inl1_inl2_inl1);
  assign c1700 = (c1693 && c576_inl2_inl1);
  assign c1701 = (c1693 && !c576_inl2_inl1);
  assign c1702 = (c1697 && c587_inl2_inl2);
  assign c1703 = (c1697 && !c587_inl2_inl2);
  assign c1704 = (c1701 && c587_inl2_inl2_inl1);
  assign c1705 = (c1701 && !c587_inl2_inl2_inl1);
  assign c1706 = (c1695 && c597_inl1_inl2);
  assign c1707 = (c1699 && c597_inl1_inl2_inl1);
  assign c1708 = (c1706 && c599_inl1_inl2);
  assign c1709 = (c1706 && !c599_inl1_inl2);
  assign c1710 = (c1703 && c597_inl2_inl2);
  assign c1711 = (c1707 && c599_inl1_inl2_inl1);
  assign c1712 = (c1707 && !c599_inl1_inl2_inl1);
  assign c1713 = (c1705 && c597_inl2_inl2_inl1);
  assign c1714 = (c1695 && !c597_inl1_inl2);
  assign c1715 = (c1710 && c599_inl2_inl2);
  assign c1716 = (c1710 && !c599_inl2_inl2);
  assign c1717 = (c1699 && !c597_inl1_inl2_inl1);
  assign c1718 = (c1713 && c599_inl2_inl2_inl1);
  assign c1719 = (c1713 && !c599_inl2_inl2_inl1);
  assign c1720 = (c1703 && !c597_inl2_inl2);
  assign c1721 = (c1705 && !c597_inl2_inl2_inl1);
  assign c1722 = ((c1694 || c1714) || c1708);
  assign c1723 = ((c1702 || c1720) || c1715);
  assign c1724 = ((c1698 || c1717) || c1711);
  assign c1725 = ((c1704 || c1721) || c1718);
  assign c558_inl2 = (t612 == 0);
  assign c558_inl2_inl1 = (mul_result1_inl16 == 0);
  assign c559_inl2 = (t613 == 0);
  assign c559_inl2_inl1 = (t609 == 0);
  assign c566_inl2 = (x_e_inl22 < b_e_inl22);
  assign c566_inl2_inl1 = (x_e_inl2_inl13 < b_e_inl2_inl13);
  assign c567_inl2 = (d_inl2 > 8);
  assign c567_inl2_inl1 = (d_inl2_inl1 > 8);
  assign c568_inl2 = (d_inl2 == 0);
  assign c568_inl2_inl1 = (d_inl2_inl1 == 0);
  assign c576_inl2 = (new_b_n_inl2 == 0);
  assign c576_inl2_inl1 = (new_b_n_inl2_inl1 == 0);
  assign c581_inl1_inl2 = (x_sign_inl24 == 0);
  assign c581_inl1_inl2_inl1 = (x_sign_inl2_inl15 == 0);
  assign c581_inl2_inl2 = (x_sign_inl24 == 0);
  assign c581_inl2_inl2_inl1 = (x_sign_inl2_inl15 == 0);
  assign c582_inl1_inl2 = (b_sign_inl24 == 0);
  assign c582_inl1_inl2_inl1 = (b_sign_inl2_inl15 == 0);
  assign c582_inl2_inl2 = (b_sign_inl24 == 0);
  assign c582_inl2_inl2_inl1 = (b_sign_inl2_inl15 == 0);
  assign c583_inl1_inl2 = (c581_inl1_inl2 && c582_inl1_inl2);
  assign c583_inl1_inl2_inl1 = (c581_inl1_inl2_inl1 && c582_inl1_inl2_inl1);
  assign c583_inl2_inl2 = (c581_inl2_inl2 && c582_inl2_inl2);
  assign c583_inl2_inl2_inl1 = (c581_inl2_inl2_inl1 && c582_inl2_inl2_inl1);
  assign c584_inl1_inl2 = (x_sign_inl24 == 1);
  assign c584_inl1_inl2_inl1 = (x_sign_inl2_inl15 == 1);
  assign c584_inl2_inl2 = (x_sign_inl24 == 1);
  assign c584_inl2_inl2_inl1 = (x_sign_inl2_inl15 == 1);
  assign c585_inl1_inl2 = (b_sign_inl24 == 1);
  assign c585_inl1_inl2_inl1 = (b_sign_inl2_inl15 == 1);
  assign c585_inl2_inl2 = (b_sign_inl24 == 1);
  assign c585_inl2_inl2_inl1 = (b_sign_inl2_inl15 == 1);
  assign c586_inl1_inl2 = (c584_inl1_inl2 && c585_inl1_inl2);
  assign c586_inl1_inl2_inl1 = (c584_inl1_inl2_inl1 && c585_inl1_inl2_inl1);
  assign c586_inl2_inl2 = (c584_inl2_inl2 && c585_inl2_inl2);
  assign c586_inl2_inl2_inl1 = (c584_inl2_inl2_inl1 && c585_inl2_inl2_inl1);
  assign c587_inl1_inl2 = (c583_inl1_inl2 || c586_inl1_inl2);
  assign c587_inl1_inl2_inl1 = (c583_inl1_inl2_inl1 || c586_inl1_inl2_inl1);
  assign c587_inl2_inl2 = (c583_inl2_inl2 || c586_inl2_inl2);
  assign c587_inl2_inl2_inl1 = (c583_inl2_inl2_inl1 || c586_inl2_inl2_inl1);
  assign c588_inl1_inl2 = (t569_inl2 < t570_inl2);
  assign c588_inl1_inl2_inl1 = (t569_inl2_inl1 < t570_inl2_inl1);
  assign c588_inl2_inl2 = (t577_inl2 < new_b_n_inl2);
  assign c588_inl2_inl2_inl1 = (t577_inl2_inl1 < new_b_n_inl2_inl1);
  assign c591_inl1_inl2 = (t590_inl1_inl2 != 0);
  assign c591_inl1_inl2_inl1 = (t590_inl1_inl2_inl1 != 0);
  assign c591_inl2_inl2 = (t590_inl2_inl2 != 0);
  assign c591_inl2_inl2_inl1 = (t590_inl2_inl2_inl1 != 0);
  assign c597_inl1_inl2 = (i_inl1_inl23 < 7);
  assign c597_inl1_inl2_inl1 = (i_inl1_inl2_inl14 < 7);
  assign c597_inl2_inl2 = (i_inl2_inl23 < 7);
  assign c597_inl2_inl2_inl1 = (i_inl2_inl2_inl14 < 7);
  assign c599_inl1_inl2 = (t598_inl1_inl2 != 0);
  assign c599_inl1_inl2_inl1 = (t598_inl1_inl2_inl1 != 0);
  assign c599_inl2_inl2 = (t598_inl2_inl2 != 0);
  assign c599_inl2_inl2_inl1 = (t598_inl2_inl2_inl1 != 0);
  assign c605 = (i2 < lst_len);
  assign c606 = (j3 < 10);
  assign c611 = (j6 < 10);
  assign c615_inl1_inl1 = (x == 0);
  assign c616_inl1_inl1 = (t608 == 0);
  assign c625_inl1_inl1 = (t624_inl1_inl1 != 0);
  assign c643_inl1_inl2 = (!c587_inl1_inl2 && c588_inl1_inl2);
  assign c643_inl1_inl2_inl1 = (!c587_inl1_inl2_inl1 && c588_inl1_inl2_inl1);
  assign c643_inl2_inl2 = (!c587_inl2_inl2 && c588_inl2_inl2);
  assign c643_inl2_inl2_inl1 = (!c587_inl2_inl2_inl1 && c588_inl2_inl2_inl1);
  assign c644_inl1_inl2 = (!c587_inl1_inl2 && !c588_inl1_inl2);
  assign c644_inl1_inl2_inl1 = (!c587_inl1_inl2_inl1 && !c588_inl1_inl2_inl1);
  assign c644_inl2_inl2 = (!c587_inl2_inl2 && !c588_inl2_inl2);
  assign c644_inl2_inl2_inl1 = (!c587_inl2_inl2_inl1 && !c588_inl2_inl2_inl1);
  assign d_inl2 = (x_e_inl24 - b_e_inl24);
  assign d_inl2_inl1 = (x_e_inl2_inl15 - b_e_inl2_inl15);
  assign e_inl1_inl13 = (t621_inl1_inl1 + 127);
  assign e_inl1_inl14 = (e_inl1_inl13 + 1);
  assign e_inl1_inl15 = c1204 ? e_inl1_inl14 : c1205 ? e_inl1_inl13 : 'bz;
  assign e_inl1_inl2 = x_e_inl24;
  assign e_inl1_inl2_inl1 = x_e_inl2_inl15;
  assign e_inl2_inl2 = x_e_inl24;
  assign e_inl2_inl2_inl1 = x_e_inl2_inl15;
  function [31:0] B_PARAM (
    input [31:0] B_PARAM_in
  );
  begin
    case (B_PARAM_in)
      0: begin
        B_PARAM = 49067;
      end
      1: begin
        B_PARAM = 16313;
      end
      2: begin
        B_PARAM = 16053;
      end
      3: begin
        B_PARAM = 48930;
      end
      4: begin
        B_PARAM = 15985;
      end
      5: begin
        B_PARAM = 16444;
      end
      6: begin
        B_PARAM = 48910;
      end
      7: begin
        B_PARAM = 16342;
      end
      8: begin
        B_PARAM = 49240;
      end
      9: begin
        B_PARAM = 48958;
      end
    endcase
  end
  endfunction
  function [31:0] W_PARAM (
    input [31:0] W_PARAM_in
  );
  begin
    case (W_PARAM_in)
      0: begin
        W_PARAM = 0;
      end
      1: begin
        W_PARAM = 0;
      end
      2: begin
        W_PARAM = 0;
      end
      3: begin
        W_PARAM = 0;
      end
      4: begin
        W_PARAM = 0;
      end
      5: begin
        W_PARAM = 0;
      end
      6: begin
        W_PARAM = 0;
      end
      7: begin
        W_PARAM = 0;
      end
      8: begin
        W_PARAM = 0;
      end
      9: begin
        W_PARAM = 0;
      end
      10: begin
        W_PARAM = 0;
      end
      11: begin
        W_PARAM = 0;
      end
      12: begin
        W_PARAM = 0;
      end
      13: begin
        W_PARAM = 0;
      end
      14: begin
        W_PARAM = 0;
      end
      15: begin
        W_PARAM = 0;
      end
      16: begin
        W_PARAM = 0;
      end
      17: begin
        W_PARAM = 0;
      end
      18: begin
        W_PARAM = 0;
      end
      19: begin
        W_PARAM = 0;
      end
      20: begin
        W_PARAM = 0;
      end
      21: begin
        W_PARAM = 0;
      end
      22: begin
        W_PARAM = 0;
      end
      23: begin
        W_PARAM = 0;
      end
      24: begin
        W_PARAM = 0;
      end
      25: begin
        W_PARAM = 0;
      end
      26: begin
        W_PARAM = 0;
      end
      27: begin
        W_PARAM = 0;
      end
      28: begin
        W_PARAM = 0;
      end
      29: begin
        W_PARAM = 0;
      end
      30: begin
        W_PARAM = 0;
      end
      31: begin
        W_PARAM = 0;
      end
      32: begin
        W_PARAM = 0;
      end
      33: begin
        W_PARAM = 0;
      end
      34: begin
        W_PARAM = 0;
      end
      35: begin
        W_PARAM = 0;
      end
      36: begin
        W_PARAM = 0;
      end
      37: begin
        W_PARAM = 0;
      end
      38: begin
        W_PARAM = 0;
      end
      39: begin
        W_PARAM = 0;
      end
      40: begin
        W_PARAM = 0;
      end
      41: begin
        W_PARAM = 0;
      end
      42: begin
        W_PARAM = 0;
      end
      43: begin
        W_PARAM = 0;
      end
      44: begin
        W_PARAM = 0;
      end
      45: begin
        W_PARAM = 0;
      end
      46: begin
        W_PARAM = 0;
      end
      47: begin
        W_PARAM = 0;
      end
      48: begin
        W_PARAM = 0;
      end
      49: begin
        W_PARAM = 0;
      end
      50: begin
        W_PARAM = 0;
      end
      51: begin
        W_PARAM = 0;
      end
      52: begin
        W_PARAM = 0;
      end
      53: begin
        W_PARAM = 0;
      end
      54: begin
        W_PARAM = 0;
      end
      55: begin
        W_PARAM = 0;
      end
      56: begin
        W_PARAM = 0;
      end
      57: begin
        W_PARAM = 0;
      end
      58: begin
        W_PARAM = 0;
      end
      59: begin
        W_PARAM = 0;
      end
      60: begin
        W_PARAM = 0;
      end
      61: begin
        W_PARAM = 0;
      end
      62: begin
        W_PARAM = 0;
      end
      63: begin
        W_PARAM = 0;
      end
      64: begin
        W_PARAM = 0;
      end
      65: begin
        W_PARAM = 0;
      end
      66: begin
        W_PARAM = 0;
      end
      67: begin
        W_PARAM = 0;
      end
      68: begin
        W_PARAM = 0;
      end
      69: begin
        W_PARAM = 0;
      end
      70: begin
        W_PARAM = 0;
      end
      71: begin
        W_PARAM = 0;
      end
      72: begin
        W_PARAM = 0;
      end
      73: begin
        W_PARAM = 0;
      end
      74: begin
        W_PARAM = 0;
      end
      75: begin
        W_PARAM = 0;
      end
      76: begin
        W_PARAM = 0;
      end
      77: begin
        W_PARAM = 0;
      end
      78: begin
        W_PARAM = 0;
      end
      79: begin
        W_PARAM = 0;
      end
      80: begin
        W_PARAM = 0;
      end
      81: begin
        W_PARAM = 0;
      end
      82: begin
        W_PARAM = 0;
      end
      83: begin
        W_PARAM = 0;
      end
      84: begin
        W_PARAM = 0;
      end
      85: begin
        W_PARAM = 0;
      end
      86: begin
        W_PARAM = 0;
      end
      87: begin
        W_PARAM = 0;
      end
      88: begin
        W_PARAM = 0;
      end
      89: begin
        W_PARAM = 0;
      end
      90: begin
        W_PARAM = 0;
      end
      91: begin
        W_PARAM = 0;
      end
      92: begin
        W_PARAM = 0;
      end
      93: begin
        W_PARAM = 0;
      end
      94: begin
        W_PARAM = 0;
      end
      95: begin
        W_PARAM = 0;
      end
      96: begin
        W_PARAM = 0;
      end
      97: begin
        W_PARAM = 0;
      end
      98: begin
        W_PARAM = 0;
      end
      99: begin
        W_PARAM = 0;
      end
      100: begin
        W_PARAM = 0;
      end
      101: begin
        W_PARAM = 0;
      end
      102: begin
        W_PARAM = 0;
      end
      103: begin
        W_PARAM = 0;
      end
      104: begin
        W_PARAM = 0;
      end
      105: begin
        W_PARAM = 0;
      end
      106: begin
        W_PARAM = 0;
      end
      107: begin
        W_PARAM = 0;
      end
      108: begin
        W_PARAM = 0;
      end
      109: begin
        W_PARAM = 0;
      end
      110: begin
        W_PARAM = 0;
      end
      111: begin
        W_PARAM = 0;
      end
      112: begin
        W_PARAM = 0;
      end
      113: begin
        W_PARAM = 0;
      end
      114: begin
        W_PARAM = 0;
      end
      115: begin
        W_PARAM = 0;
      end
      116: begin
        W_PARAM = 0;
      end
      117: begin
        W_PARAM = 0;
      end
      118: begin
        W_PARAM = 0;
      end
      119: begin
        W_PARAM = 0;
      end
      120: begin
        W_PARAM = 46358;
      end
      121: begin
        W_PARAM = 46387;
      end
      122: begin
        W_PARAM = 47711;
      end
      123: begin
        W_PARAM = 47185;
      end
      124: begin
        W_PARAM = 48013;
      end
      125: begin
        W_PARAM = 47250;
      end
      126: begin
        W_PARAM = 15304;
      end
      127: begin
        W_PARAM = 46174;
      end
      128: begin
        W_PARAM = 47397;
      end
      129: begin
        W_PARAM = 47660;
      end
      130: begin
        W_PARAM = 46864;
      end
      131: begin
        W_PARAM = 46534;
      end
      132: begin
        W_PARAM = 47851;
      end
      133: begin
        W_PARAM = 47343;
      end
      134: begin
        W_PARAM = 48155;
      end
      135: begin
        W_PARAM = 47392;
      end
      136: begin
        W_PARAM = 15450;
      end
      137: begin
        W_PARAM = 46338;
      end
      138: begin
        W_PARAM = 47541;
      end
      139: begin
        W_PARAM = 47804;
      end
      140: begin
        W_PARAM = 46857;
      end
      141: begin
        W_PARAM = 45663;
      end
      142: begin
        W_PARAM = 14510;
      end
      143: begin
        W_PARAM = 46764;
      end
      144: begin
        W_PARAM = 46942;
      end
      145: begin
        W_PARAM = 46212;
      end
      146: begin
        W_PARAM = 47205;
      end
      147: begin
        W_PARAM = 45839;
      end
      148: begin
        W_PARAM = 46322;
      end
      149: begin
        W_PARAM = 46476;
      end
      150: begin
        W_PARAM = 46263;
      end
      151: begin
        W_PARAM = 45077;
      end
      152: begin
        W_PARAM = 13928;
      end
      153: begin
        W_PARAM = 46182;
      end
      154: begin
        W_PARAM = 46356;
      end
      155: begin
        W_PARAM = 45616;
      end
      156: begin
        W_PARAM = 46617;
      end
      157: begin
        W_PARAM = 45246;
      end
      158: begin
        W_PARAM = 45730;
      end
      159: begin
        W_PARAM = 45882;
      end
      160: begin
        W_PARAM = 0;
      end
      161: begin
        W_PARAM = 0;
      end
      162: begin
        W_PARAM = 0;
      end
      163: begin
        W_PARAM = 0;
      end
      164: begin
        W_PARAM = 0;
      end
      165: begin
        W_PARAM = 0;
      end
      166: begin
        W_PARAM = 0;
      end
      167: begin
        W_PARAM = 0;
      end
      168: begin
        W_PARAM = 0;
      end
      169: begin
        W_PARAM = 0;
      end
      170: begin
        W_PARAM = 0;
      end
      171: begin
        W_PARAM = 0;
      end
      172: begin
        W_PARAM = 0;
      end
      173: begin
        W_PARAM = 0;
      end
      174: begin
        W_PARAM = 0;
      end
      175: begin
        W_PARAM = 0;
      end
      176: begin
        W_PARAM = 0;
      end
      177: begin
        W_PARAM = 0;
      end
      178: begin
        W_PARAM = 0;
      end
      179: begin
        W_PARAM = 0;
      end
      180: begin
        W_PARAM = 0;
      end
      181: begin
        W_PARAM = 0;
      end
      182: begin
        W_PARAM = 0;
      end
      183: begin
        W_PARAM = 0;
      end
      184: begin
        W_PARAM = 0;
      end
      185: begin
        W_PARAM = 0;
      end
      186: begin
        W_PARAM = 0;
      end
      187: begin
        W_PARAM = 0;
      end
      188: begin
        W_PARAM = 0;
      end
      189: begin
        W_PARAM = 0;
      end
      190: begin
        W_PARAM = 0;
      end
      191: begin
        W_PARAM = 0;
      end
      192: begin
        W_PARAM = 0;
      end
      193: begin
        W_PARAM = 0;
      end
      194: begin
        W_PARAM = 0;
      end
      195: begin
        W_PARAM = 0;
      end
      196: begin
        W_PARAM = 0;
      end
      197: begin
        W_PARAM = 0;
      end
      198: begin
        W_PARAM = 0;
      end
      199: begin
        W_PARAM = 0;
      end
      200: begin
        W_PARAM = 0;
      end
      201: begin
        W_PARAM = 0;
      end
      202: begin
        W_PARAM = 0;
      end
      203: begin
        W_PARAM = 0;
      end
      204: begin
        W_PARAM = 0;
      end
      205: begin
        W_PARAM = 0;
      end
      206: begin
        W_PARAM = 0;
      end
      207: begin
        W_PARAM = 0;
      end
      208: begin
        W_PARAM = 0;
      end
      209: begin
        W_PARAM = 0;
      end
      210: begin
        W_PARAM = 0;
      end
      211: begin
        W_PARAM = 0;
      end
      212: begin
        W_PARAM = 0;
      end
      213: begin
        W_PARAM = 0;
      end
      214: begin
        W_PARAM = 0;
      end
      215: begin
        W_PARAM = 0;
      end
      216: begin
        W_PARAM = 0;
      end
      217: begin
        W_PARAM = 0;
      end
      218: begin
        W_PARAM = 0;
      end
      219: begin
        W_PARAM = 0;
      end
      220: begin
        W_PARAM = 0;
      end
      221: begin
        W_PARAM = 0;
      end
      222: begin
        W_PARAM = 0;
      end
      223: begin
        W_PARAM = 0;
      end
      224: begin
        W_PARAM = 0;
      end
      225: begin
        W_PARAM = 0;
      end
      226: begin
        W_PARAM = 0;
      end
      227: begin
        W_PARAM = 0;
      end
      228: begin
        W_PARAM = 0;
      end
      229: begin
        W_PARAM = 0;
      end
      230: begin
        W_PARAM = 0;
      end
      231: begin
        W_PARAM = 0;
      end
      232: begin
        W_PARAM = 0;
      end
      233: begin
        W_PARAM = 0;
      end
      234: begin
        W_PARAM = 0;
      end
      235: begin
        W_PARAM = 0;
      end
      236: begin
        W_PARAM = 0;
      end
      237: begin
        W_PARAM = 0;
      end
      238: begin
        W_PARAM = 0;
      end
      239: begin
        W_PARAM = 0;
      end
      240: begin
        W_PARAM = 0;
      end
      241: begin
        W_PARAM = 0;
      end
      242: begin
        W_PARAM = 0;
      end
      243: begin
        W_PARAM = 0;
      end
      244: begin
        W_PARAM = 0;
      end
      245: begin
        W_PARAM = 0;
      end
      246: begin
        W_PARAM = 0;
      end
      247: begin
        W_PARAM = 0;
      end
      248: begin
        W_PARAM = 0;
      end
      249: begin
        W_PARAM = 0;
      end
      250: begin
        W_PARAM = 0;
      end
      251: begin
        W_PARAM = 0;
      end
      252: begin
        W_PARAM = 0;
      end
      253: begin
        W_PARAM = 0;
      end
      254: begin
        W_PARAM = 0;
      end
      255: begin
        W_PARAM = 0;
      end
      256: begin
        W_PARAM = 0;
      end
      257: begin
        W_PARAM = 0;
      end
      258: begin
        W_PARAM = 0;
      end
      259: begin
        W_PARAM = 0;
      end
      260: begin
        W_PARAM = 0;
      end
      261: begin
        W_PARAM = 0;
      end
      262: begin
        W_PARAM = 0;
      end
      263: begin
        W_PARAM = 0;
      end
      264: begin
        W_PARAM = 0;
      end
      265: begin
        W_PARAM = 0;
      end
      266: begin
        W_PARAM = 0;
      end
      267: begin
        W_PARAM = 0;
      end
      268: begin
        W_PARAM = 0;
      end
      269: begin
        W_PARAM = 0;
      end
      270: begin
        W_PARAM = 0;
      end
      271: begin
        W_PARAM = 0;
      end
      272: begin
        W_PARAM = 0;
      end
      273: begin
        W_PARAM = 0;
      end
      274: begin
        W_PARAM = 0;
      end
      275: begin
        W_PARAM = 0;
      end
      276: begin
        W_PARAM = 0;
      end
      277: begin
        W_PARAM = 0;
      end
      278: begin
        W_PARAM = 0;
      end
      279: begin
        W_PARAM = 0;
      end
      280: begin
        W_PARAM = 0;
      end
      281: begin
        W_PARAM = 0;
      end
      282: begin
        W_PARAM = 0;
      end
      283: begin
        W_PARAM = 0;
      end
      284: begin
        W_PARAM = 0;
      end
      285: begin
        W_PARAM = 0;
      end
      286: begin
        W_PARAM = 0;
      end
      287: begin
        W_PARAM = 0;
      end
      288: begin
        W_PARAM = 0;
      end
      289: begin
        W_PARAM = 0;
      end
      290: begin
        W_PARAM = 0;
      end
      291: begin
        W_PARAM = 0;
      end
      292: begin
        W_PARAM = 0;
      end
      293: begin
        W_PARAM = 0;
      end
      294: begin
        W_PARAM = 0;
      end
      295: begin
        W_PARAM = 0;
      end
      296: begin
        W_PARAM = 0;
      end
      297: begin
        W_PARAM = 0;
      end
      298: begin
        W_PARAM = 0;
      end
      299: begin
        W_PARAM = 0;
      end
      300: begin
        W_PARAM = 0;
      end
      301: begin
        W_PARAM = 0;
      end
      302: begin
        W_PARAM = 0;
      end
      303: begin
        W_PARAM = 0;
      end
      304: begin
        W_PARAM = 0;
      end
      305: begin
        W_PARAM = 0;
      end
      306: begin
        W_PARAM = 0;
      end
      307: begin
        W_PARAM = 0;
      end
      308: begin
        W_PARAM = 0;
      end
      309: begin
        W_PARAM = 0;
      end
      310: begin
        W_PARAM = 0;
      end
      311: begin
        W_PARAM = 0;
      end
      312: begin
        W_PARAM = 0;
      end
      313: begin
        W_PARAM = 0;
      end
      314: begin
        W_PARAM = 0;
      end
      315: begin
        W_PARAM = 0;
      end
      316: begin
        W_PARAM = 0;
      end
      317: begin
        W_PARAM = 0;
      end
      318: begin
        W_PARAM = 0;
      end
      319: begin
        W_PARAM = 0;
      end
      320: begin
        W_PARAM = 45187;
      end
      321: begin
        W_PARAM = 45724;
      end
      322: begin
        W_PARAM = 46950;
      end
      323: begin
        W_PARAM = 45217;
      end
      324: begin
        W_PARAM = 47274;
      end
      325: begin
        W_PARAM = 45680;
      end
      326: begin
        W_PARAM = 14537;
      end
      327: begin
        W_PARAM = 45842;
      end
      328: begin
        W_PARAM = 46246;
      end
      329: begin
        W_PARAM = 46402;
      end
      330: begin
        W_PARAM = 45522;
      end
      331: begin
        W_PARAM = 45925;
      end
      332: begin
        W_PARAM = 47160;
      end
      333: begin
        W_PARAM = 45432;
      end
      334: begin
        W_PARAM = 47876;
      end
      335: begin
        W_PARAM = 45873;
      end
      336: begin
        W_PARAM = 15111;
      end
      337: begin
        W_PARAM = 46384;
      end
      338: begin
        W_PARAM = 46452;
      end
      339: begin
        W_PARAM = 46611;
      end
      340: begin
        W_PARAM = 46303;
      end
      341: begin
        W_PARAM = 45001;
      end
      342: begin
        W_PARAM = 47600;
      end
      343: begin
        W_PARAM = 46639;
      end
      344: begin
        W_PARAM = 48693;
      end
      345: begin
        W_PARAM = 46854;
      end
      346: begin
        W_PARAM = 15925;
      end
      347: begin
        W_PARAM = 47106;
      end
      348: begin
        W_PARAM = 46074;
      end
      349: begin
        W_PARAM = 47132;
      end
      350: begin
        W_PARAM = 46836;
      end
      351: begin
        W_PARAM = 47364;
      end
      352: begin
        W_PARAM = 47778;
      end
      353: begin
        W_PARAM = 46838;
      end
      354: begin
        W_PARAM = 48825;
      end
      355: begin
        W_PARAM = 46945;
      end
      356: begin
        W_PARAM = 16058;
      end
      357: begin
        W_PARAM = 47818;
      end
      358: begin
        W_PARAM = 47190;
      end
      359: begin
        W_PARAM = 47496;
      end
      360: begin
        W_PARAM = 47170;
      end
      361: begin
        W_PARAM = 48072;
      end
      362: begin
        W_PARAM = 47781;
      end
      363: begin
        W_PARAM = 47406;
      end
      364: begin
        W_PARAM = 48842;
      end
      365: begin
        W_PARAM = 47231;
      end
      366: begin
        W_PARAM = 16085;
      end
      367: begin
        W_PARAM = 48169;
      end
      368: begin
        W_PARAM = 47723;
      end
      369: begin
        W_PARAM = 47974;
      end
      370: begin
        W_PARAM = 47403;
      end
      371: begin
        W_PARAM = 48028;
      end
      372: begin
        W_PARAM = 48019;
      end
      373: begin
        W_PARAM = 47314;
      end
      374: begin
        W_PARAM = 48655;
      end
      375: begin
        W_PARAM = 47506;
      end
      376: begin
        W_PARAM = 15912;
      end
      377: begin
        W_PARAM = 47961;
      end
      378: begin
        W_PARAM = 47723;
      end
      379: begin
        W_PARAM = 48172;
      end
      380: begin
        W_PARAM = 47938;
      end
      381: begin
        W_PARAM = 47900;
      end
      382: begin
        W_PARAM = 48319;
      end
      383: begin
        W_PARAM = 47404;
      end
      384: begin
        W_PARAM = 48604;
      end
      385: begin
        W_PARAM = 47786;
      end
      386: begin
        W_PARAM = 15898;
      end
      387: begin
        W_PARAM = 47684;
      end
      388: begin
        W_PARAM = 47607;
      end
      389: begin
        W_PARAM = 48187;
      end
      390: begin
        W_PARAM = 15884;
      end
      391: begin
        W_PARAM = 47375;
      end
      392: begin
        W_PARAM = 48603;
      end
      393: begin
        W_PARAM = 47525;
      end
      394: begin
        W_PARAM = 48745;
      end
      395: begin
        W_PARAM = 47778;
      end
      396: begin
        W_PARAM = 16008;
      end
      397: begin
        W_PARAM = 48367;
      end
      398: begin
        W_PARAM = 47786;
      end
      399: begin
        W_PARAM = 48401;
      end
      400: begin
        W_PARAM = 16017;
      end
      401: begin
        W_PARAM = 47686;
      end
      402: begin
        W_PARAM = 48582;
      end
      403: begin
        W_PARAM = 48053;
      end
      404: begin
        W_PARAM = 48901;
      end
      405: begin
        W_PARAM = 48275;
      end
      406: begin
        W_PARAM = 16130;
      end
      407: begin
        W_PARAM = 48558;
      end
      408: begin
        W_PARAM = 47876;
      end
      409: begin
        W_PARAM = 48515;
      end
      410: begin
        W_PARAM = 15857;
      end
      411: begin
        W_PARAM = 47668;
      end
      412: begin
        W_PARAM = 48450;
      end
      413: begin
        W_PARAM = 47880;
      end
      414: begin
        W_PARAM = 48713;
      end
      415: begin
        W_PARAM = 48260;
      end
      416: begin
        W_PARAM = 15943;
      end
      417: begin
        W_PARAM = 48340;
      end
      418: begin
        W_PARAM = 47889;
      end
      419: begin
        W_PARAM = 48302;
      end
      420: begin
        W_PARAM = 48019;
      end
      421: begin
        W_PARAM = 15660;
      end
      422: begin
        W_PARAM = 15620;
      end
      423: begin
        W_PARAM = 48170;
      end
      424: begin
        W_PARAM = 15548;
      end
      425: begin
        W_PARAM = 48152;
      end
      426: begin
        W_PARAM = 48506;
      end
      427: begin
        W_PARAM = 47749;
      end
      428: begin
        W_PARAM = 48047;
      end
      429: begin
        W_PARAM = 48060;
      end
      430: begin
        W_PARAM = 15864;
      end
      431: begin
        W_PARAM = 15734;
      end
      432: begin
        W_PARAM = 15911;
      end
      433: begin
        W_PARAM = 48225;
      end
      434: begin
        W_PARAM = 48849;
      end
      435: begin
        W_PARAM = 48221;
      end
      436: begin
        W_PARAM = 15899;
      end
      437: begin
        W_PARAM = 47846;
      end
      438: begin
        W_PARAM = 48023;
      end
      439: begin
        W_PARAM = 48476;
      end
      440: begin
        W_PARAM = 16047;
      end
      441: begin
        W_PARAM = 48548;
      end
      442: begin
        W_PARAM = 16037;
      end
      443: begin
        W_PARAM = 48025;
      end
      444: begin
        W_PARAM = 48868;
      end
      445: begin
        W_PARAM = 48260;
      end
      446: begin
        W_PARAM = 15609;
      end
      447: begin
        W_PARAM = 47942;
      end
      448: begin
        W_PARAM = 48068;
      end
      449: begin
        W_PARAM = 48656;
      end
      450: begin
        W_PARAM = 15912;
      end
      451: begin
        W_PARAM = 48338;
      end
      452: begin
        W_PARAM = 15688;
      end
      453: begin
        W_PARAM = 47839;
      end
      454: begin
        W_PARAM = 48686;
      end
      455: begin
        W_PARAM = 48088;
      end
      456: begin
        W_PARAM = 15764;
      end
      457: begin
        W_PARAM = 47896;
      end
      458: begin
        W_PARAM = 48127;
      end
      459: begin
        W_PARAM = 48529;
      end
      460: begin
        W_PARAM = 47754;
      end
      461: begin
        W_PARAM = 47776;
      end
      462: begin
        W_PARAM = 48481;
      end
      463: begin
        W_PARAM = 47476;
      end
      464: begin
        W_PARAM = 48404;
      end
      465: begin
        W_PARAM = 48216;
      end
      466: begin
        W_PARAM = 15846;
      end
      467: begin
        W_PARAM = 47498;
      end
      468: begin
        W_PARAM = 47955;
      end
      469: begin
        W_PARAM = 47879;
      end
      470: begin
        W_PARAM = 47600;
      end
      471: begin
        W_PARAM = 46799;
      end
      472: begin
        W_PARAM = 48418;
      end
      473: begin
        W_PARAM = 47390;
      end
      474: begin
        W_PARAM = 48685;
      end
      475: begin
        W_PARAM = 48178;
      end
      476: begin
        W_PARAM = 15973;
      end
      477: begin
        W_PARAM = 47373;
      end
      478: begin
        W_PARAM = 47865;
      end
      479: begin
        W_PARAM = 47839;
      end
      480: begin
        W_PARAM = 47425;
      end
      481: begin
        W_PARAM = 46994;
      end
      482: begin
        W_PARAM = 48255;
      end
      483: begin
        W_PARAM = 47418;
      end
      484: begin
        W_PARAM = 48666;
      end
      485: begin
        W_PARAM = 48002;
      end
      486: begin
        W_PARAM = 15927;
      end
      487: begin
        W_PARAM = 47252;
      end
      488: begin
        W_PARAM = 47936;
      end
      489: begin
        W_PARAM = 48054;
      end
      490: begin
        W_PARAM = 47252;
      end
      491: begin
        W_PARAM = 47150;
      end
      492: begin
        W_PARAM = 48029;
      end
      493: begin
        W_PARAM = 47079;
      end
      494: begin
        W_PARAM = 48591;
      end
      495: begin
        W_PARAM = 47718;
      end
      496: begin
        W_PARAM = 15839;
      end
      497: begin
        W_PARAM = 46375;
      end
      498: begin
        W_PARAM = 47745;
      end
      499: begin
        W_PARAM = 47680;
      end
      500: begin
        W_PARAM = 46881;
      end
      501: begin
        W_PARAM = 46695;
      end
      502: begin
        W_PARAM = 47566;
      end
      503: begin
        W_PARAM = 46583;
      end
      504: begin
        W_PARAM = 48689;
      end
      505: begin
        W_PARAM = 46801;
      end
      506: begin
        W_PARAM = 15922;
      end
      507: begin
        W_PARAM = 46860;
      end
      508: begin
        W_PARAM = 47323;
      end
      509: begin
        W_PARAM = 47512;
      end
      510: begin
        W_PARAM = 45781;
      end
      511: begin
        W_PARAM = 45779;
      end
      512: begin
        W_PARAM = 47492;
      end
      513: begin
        W_PARAM = 45612;
      end
      514: begin
        W_PARAM = 48594;
      end
      515: begin
        W_PARAM = 46744;
      end
      516: begin
        W_PARAM = 15828;
      end
      517: begin
        W_PARAM = 46916;
      end
      518: begin
        W_PARAM = 47139;
      end
      519: begin
        W_PARAM = 47491;
      end
      520: begin
        W_PARAM = 0;
      end
      521: begin
        W_PARAM = 0;
      end
      522: begin
        W_PARAM = 0;
      end
      523: begin
        W_PARAM = 0;
      end
      524: begin
        W_PARAM = 0;
      end
      525: begin
        W_PARAM = 0;
      end
      526: begin
        W_PARAM = 0;
      end
      527: begin
        W_PARAM = 0;
      end
      528: begin
        W_PARAM = 0;
      end
      529: begin
        W_PARAM = 0;
      end
      530: begin
        W_PARAM = 0;
      end
      531: begin
        W_PARAM = 0;
      end
      532: begin
        W_PARAM = 0;
      end
      533: begin
        W_PARAM = 0;
      end
      534: begin
        W_PARAM = 0;
      end
      535: begin
        W_PARAM = 0;
      end
      536: begin
        W_PARAM = 0;
      end
      537: begin
        W_PARAM = 0;
      end
      538: begin
        W_PARAM = 0;
      end
      539: begin
        W_PARAM = 0;
      end
      540: begin
        W_PARAM = 0;
      end
      541: begin
        W_PARAM = 0;
      end
      542: begin
        W_PARAM = 0;
      end
      543: begin
        W_PARAM = 0;
      end
      544: begin
        W_PARAM = 0;
      end
      545: begin
        W_PARAM = 0;
      end
      546: begin
        W_PARAM = 0;
      end
      547: begin
        W_PARAM = 0;
      end
      548: begin
        W_PARAM = 0;
      end
      549: begin
        W_PARAM = 0;
      end
      550: begin
        W_PARAM = 0;
      end
      551: begin
        W_PARAM = 0;
      end
      552: begin
        W_PARAM = 0;
      end
      553: begin
        W_PARAM = 0;
      end
      554: begin
        W_PARAM = 0;
      end
      555: begin
        W_PARAM = 0;
      end
      556: begin
        W_PARAM = 0;
      end
      557: begin
        W_PARAM = 0;
      end
      558: begin
        W_PARAM = 0;
      end
      559: begin
        W_PARAM = 0;
      end
      560: begin
        W_PARAM = 0;
      end
      561: begin
        W_PARAM = 0;
      end
      562: begin
        W_PARAM = 0;
      end
      563: begin
        W_PARAM = 0;
      end
      564: begin
        W_PARAM = 0;
      end
      565: begin
        W_PARAM = 0;
      end
      566: begin
        W_PARAM = 0;
      end
      567: begin
        W_PARAM = 0;
      end
      568: begin
        W_PARAM = 0;
      end
      569: begin
        W_PARAM = 0;
      end
      570: begin
        W_PARAM = 0;
      end
      571: begin
        W_PARAM = 0;
      end
      572: begin
        W_PARAM = 0;
      end
      573: begin
        W_PARAM = 0;
      end
      574: begin
        W_PARAM = 0;
      end
      575: begin
        W_PARAM = 0;
      end
      576: begin
        W_PARAM = 0;
      end
      577: begin
        W_PARAM = 0;
      end
      578: begin
        W_PARAM = 0;
      end
      579: begin
        W_PARAM = 0;
      end
      580: begin
        W_PARAM = 45709;
      end
      581: begin
        W_PARAM = 44907;
      end
      582: begin
        W_PARAM = 46479;
      end
      583: begin
        W_PARAM = 44890;
      end
      584: begin
        W_PARAM = 46762;
      end
      585: begin
        W_PARAM = 46347;
      end
      586: begin
        W_PARAM = 14291;
      end
      587: begin
        W_PARAM = 43085;
      end
      588: begin
        W_PARAM = 47002;
      end
      589: begin
        W_PARAM = 46007;
      end
      590: begin
        W_PARAM = 15542;
      end
      591: begin
        W_PARAM = 44502;
      end
      592: begin
        W_PARAM = 47075;
      end
      593: begin
        W_PARAM = 46419;
      end
      594: begin
        W_PARAM = 48300;
      end
      595: begin
        W_PARAM = 47670;
      end
      596: begin
        W_PARAM = 15075;
      end
      597: begin
        W_PARAM = 47822;
      end
      598: begin
        W_PARAM = 46658;
      end
      599: begin
        W_PARAM = 47666;
      end
      600: begin
        W_PARAM = 15364;
      end
      601: begin
        W_PARAM = 46636;
      end
      602: begin
        W_PARAM = 47870;
      end
      603: begin
        W_PARAM = 46341;
      end
      604: begin
        W_PARAM = 48147;
      end
      605: begin
        W_PARAM = 47063;
      end
      606: begin
        W_PARAM = 15217;
      end
      607: begin
        W_PARAM = 47631;
      end
      608: begin
        W_PARAM = 47011;
      end
      609: begin
        W_PARAM = 47486;
      end
      610: begin
        W_PARAM = 47780;
      end
      611: begin
        W_PARAM = 46882;
      end
      612: begin
        W_PARAM = 14684;
      end
      613: begin
        W_PARAM = 47657;
      end
      614: begin
        W_PARAM = 48091;
      end
      615: begin
        W_PARAM = 47033;
      end
      616: begin
        W_PARAM = 15371;
      end
      617: begin
        W_PARAM = 46616;
      end
      618: begin
        W_PARAM = 47244;
      end
      619: begin
        W_PARAM = 46774;
      end
      620: begin
        W_PARAM = 48593;
      end
      621: begin
        W_PARAM = 47178;
      end
      622: begin
        W_PARAM = 47177;
      end
      623: begin
        W_PARAM = 47967;
      end
      624: begin
        W_PARAM = 48694;
      end
      625: begin
        W_PARAM = 47050;
      end
      626: begin
        W_PARAM = 16017;
      end
      627: begin
        W_PARAM = 47496;
      end
      628: begin
        W_PARAM = 47562;
      end
      629: begin
        W_PARAM = 47191;
      end
      630: begin
        W_PARAM = 48616;
      end
      631: begin
        W_PARAM = 47959;
      end
      632: begin
        W_PARAM = 48299;
      end
      633: begin
        W_PARAM = 48072;
      end
      634: begin
        W_PARAM = 48902;
      end
      635: begin
        W_PARAM = 47653;
      end
      636: begin
        W_PARAM = 16172;
      end
      637: begin
        W_PARAM = 47936;
      end
      638: begin
        W_PARAM = 47684;
      end
      639: begin
        W_PARAM = 47639;
      end
      640: begin
        W_PARAM = 48526;
      end
      641: begin
        W_PARAM = 48633;
      end
      642: begin
        W_PARAM = 15917;
      end
      643: begin
        W_PARAM = 48478;
      end
      644: begin
        W_PARAM = 48931;
      end
      645: begin
        W_PARAM = 48009;
      end
      646: begin
        W_PARAM = 16190;
      end
      647: begin
        W_PARAM = 48188;
      end
      648: begin
        W_PARAM = 48025;
      end
      649: begin
        W_PARAM = 48072;
      end
      650: begin
        W_PARAM = 48488;
      end
      651: begin
        W_PARAM = 48771;
      end
      652: begin
        W_PARAM = 16169;
      end
      653: begin
        W_PARAM = 48556;
      end
      654: begin
        W_PARAM = 48894;
      end
      655: begin
        W_PARAM = 48397;
      end
      656: begin
        W_PARAM = 16035;
      end
      657: begin
        W_PARAM = 48194;
      end
      658: begin
        W_PARAM = 48315;
      end
      659: begin
        W_PARAM = 48260;
      end
      660: begin
        W_PARAM = 48425;
      end
      661: begin
        W_PARAM = 48667;
      end
      662: begin
        W_PARAM = 16040;
      end
      663: begin
        W_PARAM = 48381;
      end
      664: begin
        W_PARAM = 48971;
      end
      665: begin
        W_PARAM = 48708;
      end
      666: begin
        W_PARAM = 16255;
      end
      667: begin
        W_PARAM = 48357;
      end
      668: begin
        W_PARAM = 48462;
      end
      669: begin
        W_PARAM = 48418;
      end
      670: begin
        W_PARAM = 48624;
      end
      671: begin
        W_PARAM = 48727;
      end
      672: begin
        W_PARAM = 16149;
      end
      673: begin
        W_PARAM = 15932;
      end
      674: begin
        W_PARAM = 48937;
      end
      675: begin
        W_PARAM = 48858;
      end
      676: begin
        W_PARAM = 16232;
      end
      677: begin
        W_PARAM = 48552;
      end
      678: begin
        W_PARAM = 48619;
      end
      679: begin
        W_PARAM = 48497;
      end
      680: begin
        W_PARAM = 48654;
      end
      681: begin
        W_PARAM = 48307;
      end
      682: begin
        W_PARAM = 16085;
      end
      683: begin
        W_PARAM = 16032;
      end
      684: begin
        W_PARAM = 49005;
      end
      685: begin
        W_PARAM = 48821;
      end
      686: begin
        W_PARAM = 16257;
      end
      687: begin
        W_PARAM = 48608;
      end
      688: begin
        W_PARAM = 48602;
      end
      689: begin
        W_PARAM = 48544;
      end
      690: begin
        W_PARAM = 48769;
      end
      691: begin
        W_PARAM = 16171;
      end
      692: begin
        W_PARAM = 48321;
      end
      693: begin
        W_PARAM = 15809;
      end
      694: begin
        W_PARAM = 48878;
      end
      695: begin
        W_PARAM = 48800;
      end
      696: begin
        W_PARAM = 16138;
      end
      697: begin
        W_PARAM = 48426;
      end
      698: begin
        W_PARAM = 48668;
      end
      699: begin
        W_PARAM = 48496;
      end
      700: begin
        W_PARAM = 48859;
      end
      701: begin
        W_PARAM = 16070;
      end
      702: begin
        W_PARAM = 15902;
      end
      703: begin
        W_PARAM = 15646;
      end
      704: begin
        W_PARAM = 48661;
      end
      705: begin
        W_PARAM = 48815;
      end
      706: begin
        W_PARAM = 16145;
      end
      707: begin
        W_PARAM = 48444;
      end
      708: begin
        W_PARAM = 48649;
      end
      709: begin
        W_PARAM = 48468;
      end
      710: begin
        W_PARAM = 48897;
      end
      711: begin
        W_PARAM = 16200;
      end
      712: begin
        W_PARAM = 16139;
      end
      713: begin
        W_PARAM = 48712;
      end
      714: begin
        W_PARAM = 48857;
      end
      715: begin
        W_PARAM = 48624;
      end
      716: begin
        W_PARAM = 15969;
      end
      717: begin
        W_PARAM = 48551;
      end
      718: begin
        W_PARAM = 48678;
      end
      719: begin
        W_PARAM = 48505;
      end
      720: begin
        W_PARAM = 48824;
      end
      721: begin
        W_PARAM = 16153;
      end
      722: begin
        W_PARAM = 16040;
      end
      723: begin
        W_PARAM = 48665;
      end
      724: begin
        W_PARAM = 48950;
      end
      725: begin
        W_PARAM = 15898;
      end
      726: begin
        W_PARAM = 16137;
      end
      727: begin
        W_PARAM = 48483;
      end
      728: begin
        W_PARAM = 48763;
      end
      729: begin
        W_PARAM = 48577;
      end
      730: begin
        W_PARAM = 48775;
      end
      731: begin
        W_PARAM = 15982;
      end
      732: begin
        W_PARAM = 48642;
      end
      733: begin
        W_PARAM = 48735;
      end
      734: begin
        W_PARAM = 48797;
      end
      735: begin
        W_PARAM = 16092;
      end
      736: begin
        W_PARAM = 16136;
      end
      737: begin
        W_PARAM = 48321;
      end
      738: begin
        W_PARAM = 48721;
      end
      739: begin
        W_PARAM = 48467;
      end
      740: begin
        W_PARAM = 48666;
      end
      741: begin
        W_PARAM = 48305;
      end
      742: begin
        W_PARAM = 15623;
      end
      743: begin
        W_PARAM = 48798;
      end
      744: begin
        W_PARAM = 48841;
      end
      745: begin
        W_PARAM = 16071;
      end
      746: begin
        W_PARAM = 16118;
      end
      747: begin
        W_PARAM = 48100;
      end
      748: begin
        W_PARAM = 15535;
      end
      749: begin
        W_PARAM = 48436;
      end
      750: begin
        W_PARAM = 48624;
      end
      751: begin
        W_PARAM = 16006;
      end
      752: begin
        W_PARAM = 48703;
      end
      753: begin
        W_PARAM = 48635;
      end
      754: begin
        W_PARAM = 48804;
      end
      755: begin
        W_PARAM = 15787;
      end
      756: begin
        W_PARAM = 16154;
      end
      757: begin
        W_PARAM = 48131;
      end
      758: begin
        W_PARAM = 48680;
      end
      759: begin
        W_PARAM = 48354;
      end
      760: begin
        W_PARAM = 48594;
      end
      761: begin
        W_PARAM = 15642;
      end
      762: begin
        W_PARAM = 15480;
      end
      763: begin
        W_PARAM = 48386;
      end
      764: begin
        W_PARAM = 48810;
      end
      765: begin
        W_PARAM = 48723;
      end
      766: begin
        W_PARAM = 16176;
      end
      767: begin
        W_PARAM = 47917;
      end
      768: begin
        W_PARAM = 48462;
      end
      769: begin
        W_PARAM = 48259;
      end
      770: begin
        W_PARAM = 48413;
      end
      771: begin
        W_PARAM = 48274;
      end
      772: begin
        W_PARAM = 15385;
      end
      773: begin
        W_PARAM = 48395;
      end
      774: begin
        W_PARAM = 48805;
      end
      775: begin
        W_PARAM = 48781;
      end
      776: begin
        W_PARAM = 16193;
      end
      777: begin
        W_PARAM = 47876;
      end
      778: begin
        W_PARAM = 48443;
      end
      779: begin
        W_PARAM = 48353;
      end
      780: begin
        W_PARAM = 48228;
      end
      781: begin
        W_PARAM = 48131;
      end
      782: begin
        W_PARAM = 48508;
      end
      783: begin
        W_PARAM = 48323;
      end
      784: begin
        W_PARAM = 48787;
      end
      785: begin
        W_PARAM = 48694;
      end
      786: begin
        W_PARAM = 16155;
      end
      787: begin
        W_PARAM = 47745;
      end
      788: begin
        W_PARAM = 48299;
      end
      789: begin
        W_PARAM = 48174;
      end
      790: begin
        W_PARAM = 48153;
      end
      791: begin
        W_PARAM = 48051;
      end
      792: begin
        W_PARAM = 48150;
      end
      793: begin
        W_PARAM = 48063;
      end
      794: begin
        W_PARAM = 48706;
      end
      795: begin
        W_PARAM = 48662;
      end
      796: begin
        W_PARAM = 16064;
      end
      797: begin
        W_PARAM = 47169;
      end
      798: begin
        W_PARAM = 48153;
      end
      799: begin
        W_PARAM = 47507;
      end
      800: begin
        W_PARAM = 47854;
      end
      801: begin
        W_PARAM = 47839;
      end
      802: begin
        W_PARAM = 15911;
      end
      803: begin
        W_PARAM = 47757;
      end
      804: begin
        W_PARAM = 48262;
      end
      805: begin
        W_PARAM = 48404;
      end
      806: begin
        W_PARAM = 48585;
      end
      807: begin
        W_PARAM = 46876;
      end
      808: begin
        W_PARAM = 48115;
      end
      809: begin
        W_PARAM = 46758;
      end
      810: begin
        W_PARAM = 46566;
      end
      811: begin
        W_PARAM = 46848;
      end
      812: begin
        W_PARAM = 15841;
      end
      813: begin
        W_PARAM = 46277;
      end
      814: begin
        W_PARAM = 47621;
      end
      815: begin
        W_PARAM = 47918;
      end
      816: begin
        W_PARAM = 48596;
      end
      817: begin
        W_PARAM = 44622;
      end
      818: begin
        W_PARAM = 47961;
      end
      819: begin
        W_PARAM = 46161;
      end
      820: begin
        W_PARAM = 0;
      end
      821: begin
        W_PARAM = 0;
      end
      822: begin
        W_PARAM = 0;
      end
      823: begin
        W_PARAM = 0;
      end
      824: begin
        W_PARAM = 0;
      end
      825: begin
        W_PARAM = 0;
      end
      826: begin
        W_PARAM = 0;
      end
      827: begin
        W_PARAM = 0;
      end
      828: begin
        W_PARAM = 0;
      end
      829: begin
        W_PARAM = 0;
      end
      830: begin
        W_PARAM = 0;
      end
      831: begin
        W_PARAM = 0;
      end
      832: begin
        W_PARAM = 0;
      end
      833: begin
        W_PARAM = 0;
      end
      834: begin
        W_PARAM = 0;
      end
      835: begin
        W_PARAM = 0;
      end
      836: begin
        W_PARAM = 0;
      end
      837: begin
        W_PARAM = 0;
      end
      838: begin
        W_PARAM = 0;
      end
      839: begin
        W_PARAM = 0;
      end
      840: begin
        W_PARAM = 0;
      end
      841: begin
        W_PARAM = 0;
      end
      842: begin
        W_PARAM = 0;
      end
      843: begin
        W_PARAM = 0;
      end
      844: begin
        W_PARAM = 0;
      end
      845: begin
        W_PARAM = 0;
      end
      846: begin
        W_PARAM = 0;
      end
      847: begin
        W_PARAM = 0;
      end
      848: begin
        W_PARAM = 0;
      end
      849: begin
        W_PARAM = 0;
      end
      850: begin
        W_PARAM = 0;
      end
      851: begin
        W_PARAM = 0;
      end
      852: begin
        W_PARAM = 0;
      end
      853: begin
        W_PARAM = 0;
      end
      854: begin
        W_PARAM = 0;
      end
      855: begin
        W_PARAM = 0;
      end
      856: begin
        W_PARAM = 0;
      end
      857: begin
        W_PARAM = 0;
      end
      858: begin
        W_PARAM = 0;
      end
      859: begin
        W_PARAM = 0;
      end
      860: begin
        W_PARAM = 45852;
      end
      861: begin
        W_PARAM = 15343;
      end
      862: begin
        W_PARAM = 47550;
      end
      863: begin
        W_PARAM = 47572;
      end
      864: begin
        W_PARAM = 46907;
      end
      865: begin
        W_PARAM = 46981;
      end
      866: begin
        W_PARAM = 48003;
      end
      867: begin
        W_PARAM = 45666;
      end
      868: begin
        W_PARAM = 47907;
      end
      869: begin
        W_PARAM = 46240;
      end
      870: begin
        W_PARAM = 15723;
      end
      871: begin
        W_PARAM = 15075;
      end
      872: begin
        W_PARAM = 47624;
      end
      873: begin
        W_PARAM = 47380;
      end
      874: begin
        W_PARAM = 48536;
      end
      875: begin
        W_PARAM = 14625;
      end
      876: begin
        W_PARAM = 15587;
      end
      877: begin
        W_PARAM = 48022;
      end
      878: begin
        W_PARAM = 47919;
      end
      879: begin
        W_PARAM = 48029;
      end
      880: begin
        W_PARAM = 48224;
      end
      881: begin
        W_PARAM = 47277;
      end
      882: begin
        W_PARAM = 48278;
      end
      883: begin
        W_PARAM = 48376;
      end
      884: begin
        W_PARAM = 48332;
      end
      885: begin
        W_PARAM = 15775;
      end
      886: begin
        W_PARAM = 15446;
      end
      887: begin
        W_PARAM = 47922;
      end
      888: begin
        W_PARAM = 47504;
      end
      889: begin
        W_PARAM = 47665;
      end
      890: begin
        W_PARAM = 48728;
      end
      891: begin
        W_PARAM = 48323;
      end
      892: begin
        W_PARAM = 48464;
      end
      893: begin
        W_PARAM = 16107;
      end
      894: begin
        W_PARAM = 48372;
      end
      895: begin
        W_PARAM = 48726;
      end
      896: begin
        W_PARAM = 15791;
      end
      897: begin
        W_PARAM = 47827;
      end
      898: begin
        W_PARAM = 48283;
      end
      899: begin
        W_PARAM = 47624;
      end
      900: begin
        W_PARAM = 48816;
      end
      901: begin
        W_PARAM = 48016;
      end
      902: begin
        W_PARAM = 15088;
      end
      903: begin
        W_PARAM = 16037;
      end
      904: begin
        W_PARAM = 48846;
      end
      905: begin
        W_PARAM = 48615;
      end
      906: begin
        W_PARAM = 16150;
      end
      907: begin
        W_PARAM = 48032;
      end
      908: begin
        W_PARAM = 48421;
      end
      909: begin
        W_PARAM = 47852;
      end
      910: begin
        W_PARAM = 48849;
      end
      911: begin
        W_PARAM = 48475;
      end
      912: begin
        W_PARAM = 15816;
      end
      913: begin
        W_PARAM = 16107;
      end
      914: begin
        W_PARAM = 48882;
      end
      915: begin
        W_PARAM = 48601;
      end
      916: begin
        W_PARAM = 16156;
      end
      917: begin
        W_PARAM = 48444;
      end
      918: begin
        W_PARAM = 48547;
      end
      919: begin
        W_PARAM = 47946;
      end
      920: begin
        W_PARAM = 48443;
      end
      921: begin
        W_PARAM = 48711;
      end
      922: begin
        W_PARAM = 16007;
      end
      923: begin
        W_PARAM = 16179;
      end
      924: begin
        W_PARAM = 48991;
      end
      925: begin
        W_PARAM = 48629;
      end
      926: begin
        W_PARAM = 16135;
      end
      927: begin
        W_PARAM = 48691;
      end
      928: begin
        W_PARAM = 48495;
      end
      929: begin
        W_PARAM = 48335;
      end
      930: begin
        W_PARAM = 48721;
      end
      931: begin
        W_PARAM = 48779;
      end
      932: begin
        W_PARAM = 16271;
      end
      933: begin
        W_PARAM = 15959;
      end
      934: begin
        W_PARAM = 49042;
      end
      935: begin
        W_PARAM = 48632;
      end
      936: begin
        W_PARAM = 16146;
      end
      937: begin
        W_PARAM = 48668;
      end
      938: begin
        W_PARAM = 15745;
      end
      939: begin
        W_PARAM = 48530;
      end
      940: begin
        W_PARAM = 48607;
      end
      941: begin
        W_PARAM = 48856;
      end
      942: begin
        W_PARAM = 16104;
      end
      943: begin
        W_PARAM = 16120;
      end
      944: begin
        W_PARAM = 48947;
      end
      945: begin
        W_PARAM = 15765;
      end
      946: begin
        W_PARAM = 16154;
      end
      947: begin
        W_PARAM = 48800;
      end
      948: begin
        W_PARAM = 15657;
      end
      949: begin
        W_PARAM = 48610;
      end
      950: begin
        W_PARAM = 15953;
      end
      951: begin
        W_PARAM = 48969;
      end
      952: begin
        W_PARAM = 16203;
      end
      953: begin
        W_PARAM = 16265;
      end
      954: begin
        W_PARAM = 48992;
      end
      955: begin
        W_PARAM = 48758;
      end
      956: begin
        W_PARAM = 16176;
      end
      957: begin
        W_PARAM = 48900;
      end
      958: begin
        W_PARAM = 48684;
      end
      959: begin
        W_PARAM = 48685;
      end
      960: begin
        W_PARAM = 15781;
      end
      961: begin
        W_PARAM = 48426;
      end
      962: begin
        W_PARAM = 16136;
      end
      963: begin
        W_PARAM = 16279;
      end
      964: begin
        W_PARAM = 49098;
      end
      965: begin
        W_PARAM = 15987;
      end
      966: begin
        W_PARAM = 16038;
      end
      967: begin
        W_PARAM = 48809;
      end
      968: begin
        W_PARAM = 48644;
      end
      969: begin
        W_PARAM = 48780;
      end
      970: begin
        W_PARAM = 16142;
      end
      971: begin
        W_PARAM = 15759;
      end
      972: begin
        W_PARAM = 16259;
      end
      973: begin
        W_PARAM = 16011;
      end
      974: begin
        W_PARAM = 49154;
      end
      975: begin
        W_PARAM = 15812;
      end
      976: begin
        W_PARAM = 16157;
      end
      977: begin
        W_PARAM = 48812;
      end
      978: begin
        W_PARAM = 15935;
      end
      979: begin
        W_PARAM = 48868;
      end
      980: begin
        W_PARAM = 16139;
      end
      981: begin
        W_PARAM = 48881;
      end
      982: begin
        W_PARAM = 16087;
      end
      983: begin
        W_PARAM = 16286;
      end
      984: begin
        W_PARAM = 49035;
      end
      985: begin
        W_PARAM = 15841;
      end
      986: begin
        W_PARAM = 16075;
      end
      987: begin
        W_PARAM = 48824;
      end
      988: begin
        W_PARAM = 48771;
      end
      989: begin
        W_PARAM = 48904;
      end
      990: begin
        W_PARAM = 15892;
      end
      991: begin
        W_PARAM = 15681;
      end
      992: begin
        W_PARAM = 16028;
      end
      993: begin
        W_PARAM = 16182;
      end
      994: begin
        W_PARAM = 48966;
      end
      995: begin
        W_PARAM = 16129;
      end
      996: begin
        W_PARAM = 16027;
      end
      997: begin
        W_PARAM = 48830;
      end
      998: begin
        W_PARAM = 48776;
      end
      999: begin
        W_PARAM = 48923;
      end
      1000: begin
        W_PARAM = 16035;
      end
      1001: begin
        W_PARAM = 16076;
      end
      1002: begin
        W_PARAM = 16080;
      end
      1003: begin
        W_PARAM = 16142;
      end
      1004: begin
        W_PARAM = 48985;
      end
      1005: begin
        W_PARAM = 48623;
      end
      1006: begin
        W_PARAM = 15848;
      end
      1007: begin
        W_PARAM = 48788;
      end
      1008: begin
        W_PARAM = 48551;
      end
      1009: begin
        W_PARAM = 48875;
      end
      1010: begin
        W_PARAM = 15858;
      end
      1011: begin
        W_PARAM = 48642;
      end
      1012: begin
        W_PARAM = 16080;
      end
      1013: begin
        W_PARAM = 16004;
      end
      1014: begin
        W_PARAM = 48898;
      end
      1015: begin
        W_PARAM = 16001;
      end
      1016: begin
        W_PARAM = 48581;
      end
      1017: begin
        W_PARAM = 48645;
      end
      1018: begin
        W_PARAM = 15746;
      end
      1019: begin
        W_PARAM = 48754;
      end
      1020: begin
        W_PARAM = 48689;
      end
      1021: begin
        W_PARAM = 48919;
      end
      1022: begin
        W_PARAM = 48826;
      end
      1023: begin
        W_PARAM = 16176;
      end
      1024: begin
        W_PARAM = 48929;
      end
      1025: begin
        W_PARAM = 16075;
      end
      1026: begin
        W_PARAM = 15995;
      end
      1027: begin
        W_PARAM = 48575;
      end
      1028: begin
        W_PARAM = 16117;
      end
      1029: begin
        W_PARAM = 15656;
      end
      1030: begin
        W_PARAM = 48776;
      end
      1031: begin
        W_PARAM = 48665;
      end
      1032: begin
        W_PARAM = 48573;
      end
      1033: begin
        W_PARAM = 16146;
      end
      1034: begin
        W_PARAM = 48686;
      end
      1035: begin
        W_PARAM = 16002;
      end
      1036: begin
        W_PARAM = 16058;
      end
      1037: begin
        W_PARAM = 48462;
      end
      1038: begin
        W_PARAM = 48833;
      end
      1039: begin
        W_PARAM = 48559;
      end
      1040: begin
        W_PARAM = 48600;
      end
      1041: begin
        W_PARAM = 48842;
      end
      1042: begin
        W_PARAM = 48840;
      end
      1043: begin
        W_PARAM = 16269;
      end
      1044: begin
        W_PARAM = 48770;
      end
      1045: begin
        W_PARAM = 16135;
      end
      1046: begin
        W_PARAM = 48421;
      end
      1047: begin
        W_PARAM = 48584;
      end
      1048: begin
        W_PARAM = 48777;
      end
      1049: begin
        W_PARAM = 48542;
      end
      1050: begin
        W_PARAM = 48818;
      end
      1051: begin
        W_PARAM = 48855;
      end
      1052: begin
        W_PARAM = 48570;
      end
      1053: begin
        W_PARAM = 48837;
      end
      1054: begin
        W_PARAM = 48725;
      end
      1055: begin
        W_PARAM = 16202;
      end
      1056: begin
        W_PARAM = 16109;
      end
      1057: begin
        W_PARAM = 48527;
      end
      1058: begin
        W_PARAM = 16035;
      end
      1059: begin
        W_PARAM = 48453;
      end
      1060: begin
        W_PARAM = 48747;
      end
      1061: begin
        W_PARAM = 48821;
      end
      1062: begin
        W_PARAM = 48732;
      end
      1063: begin
        W_PARAM = 48947;
      end
      1064: begin
        W_PARAM = 15805;
      end
      1065: begin
        W_PARAM = 16032;
      end
      1066: begin
        W_PARAM = 16178;
      end
      1067: begin
        W_PARAM = 48252;
      end
      1068: begin
        W_PARAM = 16087;
      end
      1069: begin
        W_PARAM = 48127;
      end
      1070: begin
        W_PARAM = 48553;
      end
      1071: begin
        W_PARAM = 48796;
      end
      1072: begin
        W_PARAM = 48803;
      end
      1073: begin
        W_PARAM = 48856;
      end
      1074: begin
        W_PARAM = 15835;
      end
      1075: begin
        W_PARAM = 48810;
      end
      1076: begin
        W_PARAM = 16235;
      end
      1077: begin
        W_PARAM = 47867;
      end
      1078: begin
        W_PARAM = 16097;
      end
      1079: begin
        W_PARAM = 47814;
      end
      1080: begin
        W_PARAM = 48305;
      end
      1081: begin
        W_PARAM = 48784;
      end
      1082: begin
        W_PARAM = 15640;
      end
      1083: begin
        W_PARAM = 48639;
      end
      1084: begin
        W_PARAM = 48499;
      end
      1085: begin
        W_PARAM = 47902;
      end
      1086: begin
        W_PARAM = 16061;
      end
      1087: begin
        W_PARAM = 47340;
      end
      1088: begin
        W_PARAM = 15788;
      end
      1089: begin
        W_PARAM = 47534;
      end
      1090: begin
        W_PARAM = 15397;
      end
      1091: begin
        W_PARAM = 48609;
      end
      1092: begin
        W_PARAM = 15816;
      end
      1093: begin
        W_PARAM = 47399;
      end
      1094: begin
        W_PARAM = 47745;
      end
      1095: begin
        W_PARAM = 16027;
      end
      1096: begin
        W_PARAM = 48803;
      end
      1097: begin
        W_PARAM = 46485;
      end
      1098: begin
        W_PARAM = 15509;
      end
      1099: begin
        W_PARAM = 47152;
      end
      1100: begin
        W_PARAM = 47892;
      end
      1101: begin
        W_PARAM = 48662;
      end
      1102: begin
        W_PARAM = 47559;
      end
      1103: begin
        W_PARAM = 46484;
      end
      1104: begin
        W_PARAM = 47614;
      end
      1105: begin
        W_PARAM = 15699;
      end
      1106: begin
        W_PARAM = 15840;
      end
      1107: begin
        W_PARAM = 45345;
      end
      1108: begin
        W_PARAM = 48195;
      end
      1109: begin
        W_PARAM = 46084;
      end
      1110: begin
        W_PARAM = 0;
      end
      1111: begin
        W_PARAM = 0;
      end
      1112: begin
        W_PARAM = 0;
      end
      1113: begin
        W_PARAM = 0;
      end
      1114: begin
        W_PARAM = 0;
      end
      1115: begin
        W_PARAM = 0;
      end
      1116: begin
        W_PARAM = 0;
      end
      1117: begin
        W_PARAM = 0;
      end
      1118: begin
        W_PARAM = 0;
      end
      1119: begin
        W_PARAM = 0;
      end
      1120: begin
        W_PARAM = 0;
      end
      1121: begin
        W_PARAM = 0;
      end
      1122: begin
        W_PARAM = 0;
      end
      1123: begin
        W_PARAM = 0;
      end
      1124: begin
        W_PARAM = 0;
      end
      1125: begin
        W_PARAM = 0;
      end
      1126: begin
        W_PARAM = 0;
      end
      1127: begin
        W_PARAM = 0;
      end
      1128: begin
        W_PARAM = 0;
      end
      1129: begin
        W_PARAM = 0;
      end
      1130: begin
        W_PARAM = 45466;
      end
      1131: begin
        W_PARAM = 45409;
      end
      1132: begin
        W_PARAM = 47105;
      end
      1133: begin
        W_PARAM = 14446;
      end
      1134: begin
        W_PARAM = 45993;
      end
      1135: begin
        W_PARAM = 47049;
      end
      1136: begin
        W_PARAM = 45078;
      end
      1137: begin
        W_PARAM = 45045;
      end
      1138: begin
        W_PARAM = 46608;
      end
      1139: begin
        W_PARAM = 45199;
      end
      1140: begin
        W_PARAM = 47003;
      end
      1141: begin
        W_PARAM = 15565;
      end
      1142: begin
        W_PARAM = 48075;
      end
      1143: begin
        W_PARAM = 15234;
      end
      1144: begin
        W_PARAM = 46836;
      end
      1145: begin
        W_PARAM = 48084;
      end
      1146: begin
        W_PARAM = 48229;
      end
      1147: begin
        W_PARAM = 45894;
      end
      1148: begin
        W_PARAM = 47894;
      end
      1149: begin
        W_PARAM = 46472;
      end
      1150: begin
        W_PARAM = 47857;
      end
      1151: begin
        W_PARAM = 15243;
      end
      1152: begin
        W_PARAM = 48373;
      end
      1153: begin
        W_PARAM = 15781;
      end
      1154: begin
        W_PARAM = 48247;
      end
      1155: begin
        W_PARAM = 48290;
      end
      1156: begin
        W_PARAM = 48214;
      end
      1157: begin
        W_PARAM = 15149;
      end
      1158: begin
        W_PARAM = 48020;
      end
      1159: begin
        W_PARAM = 47950;
      end
      1160: begin
        W_PARAM = 48263;
      end
      1161: begin
        W_PARAM = 15635;
      end
      1162: begin
        W_PARAM = 48714;
      end
      1163: begin
        W_PARAM = 15932;
      end
      1164: begin
        W_PARAM = 15764;
      end
      1165: begin
        W_PARAM = 48667;
      end
      1166: begin
        W_PARAM = 15802;
      end
      1167: begin
        W_PARAM = 48000;
      end
      1168: begin
        W_PARAM = 48221;
      end
      1169: begin
        W_PARAM = 47661;
      end
      1170: begin
        W_PARAM = 48808;
      end
      1171: begin
        W_PARAM = 15960;
      end
      1172: begin
        W_PARAM = 15825;
      end
      1173: begin
        W_PARAM = 16212;
      end
      1174: begin
        W_PARAM = 15825;
      end
      1175: begin
        W_PARAM = 48949;
      end
      1176: begin
        W_PARAM = 15961;
      end
      1177: begin
        W_PARAM = 48773;
      end
      1178: begin
        W_PARAM = 48664;
      end
      1179: begin
        W_PARAM = 48185;
      end
      1180: begin
        W_PARAM = 48842;
      end
      1181: begin
        W_PARAM = 15987;
      end
      1182: begin
        W_PARAM = 16216;
      end
      1183: begin
        W_PARAM = 16141;
      end
      1184: begin
        W_PARAM = 48773;
      end
      1185: begin
        W_PARAM = 48904;
      end
      1186: begin
        W_PARAM = 15830;
      end
      1187: begin
        W_PARAM = 48785;
      end
      1188: begin
        W_PARAM = 48770;
      end
      1189: begin
        W_PARAM = 48223;
      end
      1190: begin
        W_PARAM = 15461;
      end
      1191: begin
        W_PARAM = 15351;
      end
      1192: begin
        W_PARAM = 15997;
      end
      1193: begin
        W_PARAM = 16057;
      end
      1194: begin
        W_PARAM = 48518;
      end
      1195: begin
        W_PARAM = 15602;
      end
      1196: begin
        W_PARAM = 48539;
      end
      1197: begin
        W_PARAM = 48794;
      end
      1198: begin
        W_PARAM = 48663;
      end
      1199: begin
        W_PARAM = 48526;
      end
      1200: begin
        W_PARAM = 15887;
      end
      1201: begin
        W_PARAM = 15928;
      end
      1202: begin
        W_PARAM = 16038;
      end
      1203: begin
        W_PARAM = 16208;
      end
      1204: begin
        W_PARAM = 48904;
      end
      1205: begin
        W_PARAM = 48933;
      end
      1206: begin
        W_PARAM = 15958;
      end
      1207: begin
        W_PARAM = 48846;
      end
      1208: begin
        W_PARAM = 15856;
      end
      1209: begin
        W_PARAM = 48721;
      end
      1210: begin
        W_PARAM = 16110;
      end
      1211: begin
        W_PARAM = 15961;
      end
      1212: begin
        W_PARAM = 16194;
      end
      1213: begin
        W_PARAM = 16053;
      end
      1214: begin
        W_PARAM = 48924;
      end
      1215: begin
        W_PARAM = 48852;
      end
      1216: begin
        W_PARAM = 48674;
      end
      1217: begin
        W_PARAM = 48949;
      end
      1218: begin
        W_PARAM = 16124;
      end
      1219: begin
        W_PARAM = 48839;
      end
      1220: begin
        W_PARAM = 15905;
      end
      1221: begin
        W_PARAM = 16033;
      end
      1222: begin
        W_PARAM = 16081;
      end
      1223: begin
        W_PARAM = 16196;
      end
      1224: begin
        W_PARAM = 48938;
      end
      1225: begin
        W_PARAM = 48181;
      end
      1226: begin
        W_PARAM = 48455;
      end
      1227: begin
        W_PARAM = 49030;
      end
      1228: begin
        W_PARAM = 16120;
      end
      1229: begin
        W_PARAM = 48822;
      end
      1230: begin
        W_PARAM = 16167;
      end
      1231: begin
        W_PARAM = 48723;
      end
      1232: begin
        W_PARAM = 16135;
      end
      1233: begin
        W_PARAM = 16177;
      end
      1234: begin
        W_PARAM = 48888;
      end
      1235: begin
        W_PARAM = 16116;
      end
      1236: begin
        W_PARAM = 48708;
      end
      1237: begin
        W_PARAM = 49030;
      end
      1238: begin
        W_PARAM = 15932;
      end
      1239: begin
        W_PARAM = 48923;
      end
      1240: begin
        W_PARAM = 48680;
      end
      1241: begin
        W_PARAM = 48663;
      end
      1242: begin
        W_PARAM = 16135;
      end
      1243: begin
        W_PARAM = 16038;
      end
      1244: begin
        W_PARAM = 48778;
      end
      1245: begin
        W_PARAM = 15903;
      end
      1246: begin
        W_PARAM = 48498;
      end
      1247: begin
        W_PARAM = 48920;
      end
      1248: begin
        W_PARAM = 16224;
      end
      1249: begin
        W_PARAM = 48934;
      end
      1250: begin
        W_PARAM = 15896;
      end
      1251: begin
        W_PARAM = 16097;
      end
      1252: begin
        W_PARAM = 15740;
      end
      1253: begin
        W_PARAM = 16135;
      end
      1254: begin
        W_PARAM = 15992;
      end
      1255: begin
        W_PARAM = 48911;
      end
      1256: begin
        W_PARAM = 15654;
      end
      1257: begin
        W_PARAM = 48912;
      end
      1258: begin
        W_PARAM = 48552;
      end
      1259: begin
        W_PARAM = 48773;
      end
      1260: begin
        W_PARAM = 48665;
      end
      1261: begin
        W_PARAM = 16042;
      end
      1262: begin
        W_PARAM = 16169;
      end
      1263: begin
        W_PARAM = 16031;
      end
      1264: begin
        W_PARAM = 48802;
      end
      1265: begin
        W_PARAM = 48606;
      end
      1266: begin
        W_PARAM = 48675;
      end
      1267: begin
        W_PARAM = 48968;
      end
      1268: begin
        W_PARAM = 16195;
      end
      1269: begin
        W_PARAM = 48908;
      end
      1270: begin
        W_PARAM = 16074;
      end
      1271: begin
        W_PARAM = 48729;
      end
      1272: begin
        W_PARAM = 15903;
      end
      1273: begin
        W_PARAM = 16065;
      end
      1274: begin
        W_PARAM = 48928;
      end
      1275: begin
        W_PARAM = 16179;
      end
      1276: begin
        W_PARAM = 48663;
      end
      1277: begin
        W_PARAM = 48957;
      end
      1278: begin
        W_PARAM = 16151;
      end
      1279: begin
        W_PARAM = 48893;
      end
      1280: begin
        W_PARAM = 48776;
      end
      1281: begin
        W_PARAM = 16024;
      end
      1282: begin
        W_PARAM = 16035;
      end
      1283: begin
        W_PARAM = 16162;
      end
      1284: begin
        W_PARAM = 48295;
      end
      1285: begin
        W_PARAM = 48433;
      end
      1286: begin
        W_PARAM = 15843;
      end
      1287: begin
        W_PARAM = 48953;
      end
      1288: begin
        W_PARAM = 16094;
      end
      1289: begin
        W_PARAM = 48957;
      end
      1290: begin
        W_PARAM = 16050;
      end
      1291: begin
        W_PARAM = 15750;
      end
      1292: begin
        W_PARAM = 15890;
      end
      1293: begin
        W_PARAM = 48060;
      end
      1294: begin
        W_PARAM = 15438;
      end
      1295: begin
        W_PARAM = 15774;
      end
      1296: begin
        W_PARAM = 15895;
      end
      1297: begin
        W_PARAM = 48935;
      end
      1298: begin
        W_PARAM = 15989;
      end
      1299: begin
        W_PARAM = 48831;
      end
      1300: begin
        W_PARAM = 15578;
      end
      1301: begin
        W_PARAM = 48912;
      end
      1302: begin
        W_PARAM = 16021;
      end
      1303: begin
        W_PARAM = 16143;
      end
      1304: begin
        W_PARAM = 48771;
      end
      1305: begin
        W_PARAM = 16206;
      end
      1306: begin
        W_PARAM = 48693;
      end
      1307: begin
        W_PARAM = 48902;
      end
      1308: begin
        W_PARAM = 15981;
      end
      1309: begin
        W_PARAM = 48845;
      end
      1310: begin
        W_PARAM = 15869;
      end
      1311: begin
        W_PARAM = 16081;
      end
      1312: begin
        W_PARAM = 48641;
      end
      1313: begin
        W_PARAM = 48501;
      end
      1314: begin
        W_PARAM = 16081;
      end
      1315: begin
        W_PARAM = 16059;
      end
      1316: begin
        W_PARAM = 48583;
      end
      1317: begin
        W_PARAM = 48786;
      end
      1318: begin
        W_PARAM = 15164;
      end
      1319: begin
        W_PARAM = 48958;
      end
      1320: begin
        W_PARAM = 15791;
      end
      1321: begin
        W_PARAM = 15617;
      end
      1322: begin
        W_PARAM = 15644;
      end
      1323: begin
        W_PARAM = 48647;
      end
      1324: begin
        W_PARAM = 16176;
      end
      1325: begin
        W_PARAM = 48936;
      end
      1326: begin
        W_PARAM = 15834;
      end
      1327: begin
        W_PARAM = 48746;
      end
      1328: begin
        W_PARAM = 16127;
      end
      1329: begin
        W_PARAM = 48860;
      end
      1330: begin
        W_PARAM = 48654;
      end
      1331: begin
        W_PARAM = 48746;
      end
      1332: begin
        W_PARAM = 48867;
      end
      1333: begin
        W_PARAM = 48821;
      end
      1334: begin
        W_PARAM = 16218;
      end
      1335: begin
        W_PARAM = 16149;
      end
      1336: begin
        W_PARAM = 16003;
      end
      1337: begin
        W_PARAM = 15635;
      end
      1338: begin
        W_PARAM = 15133;
      end
      1339: begin
        W_PARAM = 48912;
      end
      1340: begin
        W_PARAM = 15396;
      end
      1341: begin
        W_PARAM = 48852;
      end
      1342: begin
        W_PARAM = 48969;
      end
      1343: begin
        W_PARAM = 48132;
      end
      1344: begin
        W_PARAM = 16241;
      end
      1345: begin
        W_PARAM = 48650;
      end
      1346: begin
        W_PARAM = 16062;
      end
      1347: begin
        W_PARAM = 48563;
      end
      1348: begin
        W_PARAM = 16057;
      end
      1349: begin
        W_PARAM = 48771;
      end
      1350: begin
        W_PARAM = 48781;
      end
      1351: begin
        W_PARAM = 48905;
      end
      1352: begin
        W_PARAM = 48967;
      end
      1353: begin
        W_PARAM = 48975;
      end
      1354: begin
        W_PARAM = 16246;
      end
      1355: begin
        W_PARAM = 16161;
      end
      1356: begin
        W_PARAM = 16175;
      end
      1357: begin
        W_PARAM = 48380;
      end
      1358: begin
        W_PARAM = 15965;
      end
      1359: begin
        W_PARAM = 48490;
      end
      1360: begin
        W_PARAM = 48879;
      end
      1361: begin
        W_PARAM = 49026;
      end
      1362: begin
        W_PARAM = 48874;
      end
      1363: begin
        W_PARAM = 48546;
      end
      1364: begin
        W_PARAM = 16200;
      end
      1365: begin
        W_PARAM = 16286;
      end
      1366: begin
        W_PARAM = 48921;
      end
      1367: begin
        W_PARAM = 48109;
      end
      1368: begin
        W_PARAM = 16158;
      end
      1369: begin
        W_PARAM = 48223;
      end
      1370: begin
        W_PARAM = 48545;
      end
      1371: begin
        W_PARAM = 48922;
      end
      1372: begin
        W_PARAM = 15656;
      end
      1373: begin
        W_PARAM = 47989;
      end
      1374: begin
        W_PARAM = 15459;
      end
      1375: begin
        W_PARAM = 16083;
      end
      1376: begin
        W_PARAM = 48774;
      end
      1377: begin
        W_PARAM = 47851;
      end
      1378: begin
        W_PARAM = 16120;
      end
      1379: begin
        W_PARAM = 47944;
      end
      1380: begin
        W_PARAM = 48259;
      end
      1381: begin
        W_PARAM = 48564;
      end
      1382: begin
        W_PARAM = 48269;
      end
      1383: begin
        W_PARAM = 47137;
      end
      1384: begin
        W_PARAM = 48539;
      end
      1385: begin
        W_PARAM = 15809;
      end
      1386: begin
        W_PARAM = 48282;
      end
      1387: begin
        W_PARAM = 47515;
      end
      1388: begin
        W_PARAM = 15868;
      end
      1389: begin
        W_PARAM = 47781;
      end
      1390: begin
        W_PARAM = 47417;
      end
      1391: begin
        W_PARAM = 48479;
      end
      1392: begin
        W_PARAM = 48264;
      end
      1393: begin
        W_PARAM = 46778;
      end
      1394: begin
        W_PARAM = 48066;
      end
      1395: begin
        W_PARAM = 48239;
      end
      1396: begin
        W_PARAM = 15789;
      end
      1397: begin
        W_PARAM = 46929;
      end
      1398: begin
        W_PARAM = 15353;
      end
      1399: begin
        W_PARAM = 47438;
      end
      1400: begin
        W_PARAM = 0;
      end
      1401: begin
        W_PARAM = 0;
      end
      1402: begin
        W_PARAM = 0;
      end
      1403: begin
        W_PARAM = 0;
      end
      1404: begin
        W_PARAM = 0;
      end
      1405: begin
        W_PARAM = 0;
      end
      1406: begin
        W_PARAM = 0;
      end
      1407: begin
        W_PARAM = 0;
      end
      1408: begin
        W_PARAM = 0;
      end
      1409: begin
        W_PARAM = 0;
      end
      1410: begin
        W_PARAM = 0;
      end
      1411: begin
        W_PARAM = 0;
      end
      1412: begin
        W_PARAM = 0;
      end
      1413: begin
        W_PARAM = 0;
      end
      1414: begin
        W_PARAM = 0;
      end
      1415: begin
        W_PARAM = 0;
      end
      1416: begin
        W_PARAM = 0;
      end
      1417: begin
        W_PARAM = 0;
      end
      1418: begin
        W_PARAM = 0;
      end
      1419: begin
        W_PARAM = 0;
      end
      1420: begin
        W_PARAM = 47847;
      end
      1421: begin
        W_PARAM = 15191;
      end
      1422: begin
        W_PARAM = 15238;
      end
      1423: begin
        W_PARAM = 47451;
      end
      1424: begin
        W_PARAM = 47696;
      end
      1425: begin
        W_PARAM = 48001;
      end
      1426: begin
        W_PARAM = 14860;
      end
      1427: begin
        W_PARAM = 46239;
      end
      1428: begin
        W_PARAM = 47775;
      end
      1429: begin
        W_PARAM = 46271;
      end
      1430: begin
        W_PARAM = 48295;
      end
      1431: begin
        W_PARAM = 15669;
      end
      1432: begin
        W_PARAM = 48127;
      end
      1433: begin
        W_PARAM = 16056;
      end
      1434: begin
        W_PARAM = 15366;
      end
      1435: begin
        W_PARAM = 48608;
      end
      1436: begin
        W_PARAM = 48715;
      end
      1437: begin
        W_PARAM = 48311;
      end
      1438: begin
        W_PARAM = 48426;
      end
      1439: begin
        W_PARAM = 48208;
      end
      1440: begin
        W_PARAM = 48445;
      end
      1441: begin
        W_PARAM = 15829;
      end
      1442: begin
        W_PARAM = 15689;
      end
      1443: begin
        W_PARAM = 16168;
      end
      1444: begin
        W_PARAM = 15661;
      end
      1445: begin
        W_PARAM = 48930;
      end
      1446: begin
        W_PARAM = 15877;
      end
      1447: begin
        W_PARAM = 48665;
      end
      1448: begin
        W_PARAM = 48646;
      end
      1449: begin
        W_PARAM = 48293;
      end
      1450: begin
        W_PARAM = 48899;
      end
      1451: begin
        W_PARAM = 16149;
      end
      1452: begin
        W_PARAM = 15769;
      end
      1453: begin
        W_PARAM = 16231;
      end
      1454: begin
        W_PARAM = 15885;
      end
      1455: begin
        W_PARAM = 48905;
      end
      1456: begin
        W_PARAM = 48858;
      end
      1457: begin
        W_PARAM = 16042;
      end
      1458: begin
        W_PARAM = 48891;
      end
      1459: begin
        W_PARAM = 48521;
      end
      1460: begin
        W_PARAM = 15664;
      end
      1461: begin
        W_PARAM = 16095;
      end
      1462: begin
        W_PARAM = 15758;
      end
      1463: begin
        W_PARAM = 16158;
      end
      1464: begin
        W_PARAM = 48792;
      end
      1465: begin
        W_PARAM = 48923;
      end
      1466: begin
        W_PARAM = 48637;
      end
      1467: begin
        W_PARAM = 16039;
      end
      1468: begin
        W_PARAM = 48780;
      end
      1469: begin
        W_PARAM = 48706;
      end
      1470: begin
        W_PARAM = 48265;
      end
      1471: begin
        W_PARAM = 48788;
      end
      1472: begin
        W_PARAM = 15237;
      end
      1473: begin
        W_PARAM = 16143;
      end
      1474: begin
        W_PARAM = 48786;
      end
      1475: begin
        W_PARAM = 15892;
      end
      1476: begin
        W_PARAM = 48823;
      end
      1477: begin
        W_PARAM = 16007;
      end
      1478: begin
        W_PARAM = 15977;
      end
      1479: begin
        W_PARAM = 48769;
      end
      1480: begin
        W_PARAM = 15971;
      end
      1481: begin
        W_PARAM = 48949;
      end
      1482: begin
        W_PARAM = 16035;
      end
      1483: begin
        W_PARAM = 48236;
      end
      1484: begin
        W_PARAM = 47899;
      end
      1485: begin
        W_PARAM = 48774;
      end
      1486: begin
        W_PARAM = 16013;
      end
      1487: begin
        W_PARAM = 16166;
      end
      1488: begin
        W_PARAM = 48684;
      end
      1489: begin
        W_PARAM = 48798;
      end
      1490: begin
        W_PARAM = 15814;
      end
      1491: begin
        W_PARAM = 48967;
      end
      1492: begin
        W_PARAM = 48578;
      end
      1493: begin
        W_PARAM = 15971;
      end
      1494: begin
        W_PARAM = 15919;
      end
      1495: begin
        W_PARAM = 15808;
      end
      1496: begin
        W_PARAM = 15496;
      end
      1497: begin
        W_PARAM = 16132;
      end
      1498: begin
        W_PARAM = 15953;
      end
      1499: begin
        W_PARAM = 48868;
      end
      1500: begin
        W_PARAM = 16153;
      end
      1501: begin
        W_PARAM = 48811;
      end
      1502: begin
        W_PARAM = 15880;
      end
      1503: begin
        W_PARAM = 15785;
      end
      1504: begin
        W_PARAM = 48728;
      end
      1505: begin
        W_PARAM = 16030;
      end
      1506: begin
        W_PARAM = 16136;
      end
      1507: begin
        W_PARAM = 48779;
      end
      1508: begin
        W_PARAM = 48898;
      end
      1509: begin
        W_PARAM = 48806;
      end
      1510: begin
        W_PARAM = 15930;
      end
      1511: begin
        W_PARAM = 48979;
      end
      1512: begin
        W_PARAM = 16044;
      end
      1513: begin
        W_PARAM = 15811;
      end
      1514: begin
        W_PARAM = 15635;
      end
      1515: begin
        W_PARAM = 15785;
      end
      1516: begin
        W_PARAM = 48968;
      end
      1517: begin
        W_PARAM = 48812;
      end
      1518: begin
        W_PARAM = 16146;
      end
      1519: begin
        W_PARAM = 16164;
      end
      1520: begin
        W_PARAM = 48702;
      end
      1521: begin
        W_PARAM = 48945;
      end
      1522: begin
        W_PARAM = 15832;
      end
      1523: begin
        W_PARAM = 15811;
      end
      1524: begin
        W_PARAM = 16068;
      end
      1525: begin
        W_PARAM = 48623;
      end
      1526: begin
        W_PARAM = 48847;
      end
      1527: begin
        W_PARAM = 16029;
      end
      1528: begin
        W_PARAM = 16068;
      end
      1529: begin
        W_PARAM = 15863;
      end
      1530: begin
        W_PARAM = 16004;
      end
      1531: begin
        W_PARAM = 48720;
      end
      1532: begin
        W_PARAM = 15698;
      end
      1533: begin
        W_PARAM = 15895;
      end
      1534: begin
        W_PARAM = 48921;
      end
      1535: begin
        W_PARAM = 15746;
      end
      1536: begin
        W_PARAM = 48912;
      end
      1537: begin
        W_PARAM = 16036;
      end
      1538: begin
        W_PARAM = 15735;
      end
      1539: begin
        W_PARAM = 16108;
      end
      1540: begin
        W_PARAM = 15892;
      end
      1541: begin
        W_PARAM = 48771;
      end
      1542: begin
        W_PARAM = 16009;
      end
      1543: begin
        W_PARAM = 15840;
      end
      1544: begin
        W_PARAM = 15904;
      end
      1545: begin
        W_PARAM = 48733;
      end
      1546: begin
        W_PARAM = 16044;
      end
      1547: begin
        W_PARAM = 48819;
      end
      1548: begin
        W_PARAM = 16037;
      end
      1549: begin
        W_PARAM = 48900;
      end
      1550: begin
        W_PARAM = 15771;
      end
      1551: begin
        W_PARAM = 16056;
      end
      1552: begin
        W_PARAM = 15720;
      end
      1553: begin
        W_PARAM = 16004;
      end
      1554: begin
        W_PARAM = 16012;
      end
      1555: begin
        W_PARAM = 48738;
      end
      1556: begin
        W_PARAM = 48934;
      end
      1557: begin
        W_PARAM = 48933;
      end
      1558: begin
        W_PARAM = 15832;
      end
      1559: begin
        W_PARAM = 16069;
      end
      1560: begin
        W_PARAM = 15370;
      end
      1561: begin
        W_PARAM = 48831;
      end
      1562: begin
        W_PARAM = 16115;
      end
      1563: begin
        W_PARAM = 16160;
      end
      1564: begin
        W_PARAM = 15900;
      end
      1565: begin
        W_PARAM = 15831;
      end
      1566: begin
        W_PARAM = 48745;
      end
      1567: begin
        W_PARAM = 48514;
      end
      1568: begin
        W_PARAM = 15815;
      end
      1569: begin
        W_PARAM = 48972;
      end
      1570: begin
        W_PARAM = 16051;
      end
      1571: begin
        W_PARAM = 48831;
      end
      1572: begin
        W_PARAM = 15848;
      end
      1573: begin
        W_PARAM = 48674;
      end
      1574: begin
        W_PARAM = 48697;
      end
      1575: begin
        W_PARAM = 15993;
      end
      1576: begin
        W_PARAM = 48537;
      end
      1577: begin
        W_PARAM = 48795;
      end
      1578: begin
        W_PARAM = 16188;
      end
      1579: begin
        W_PARAM = 48820;
      end
      1580: begin
        W_PARAM = 16138;
      end
      1581: begin
        W_PARAM = 48709;
      end
      1582: begin
        W_PARAM = 15814;
      end
      1583: begin
        W_PARAM = 48117;
      end
      1584: begin
        W_PARAM = 15973;
      end
      1585: begin
        W_PARAM = 15881;
      end
      1586: begin
        W_PARAM = 15984;
      end
      1587: begin
        W_PARAM = 48835;
      end
      1588: begin
        W_PARAM = 48841;
      end
      1589: begin
        W_PARAM = 48771;
      end
      1590: begin
        W_PARAM = 15876;
      end
      1591: begin
        W_PARAM = 48665;
      end
      1592: begin
        W_PARAM = 48402;
      end
      1593: begin
        W_PARAM = 16016;
      end
      1594: begin
        W_PARAM = 16097;
      end
      1595: begin
        W_PARAM = 48547;
      end
      1596: begin
        W_PARAM = 16089;
      end
      1597: begin
        W_PARAM = 49013;
      end
      1598: begin
        W_PARAM = 15961;
      end
      1599: begin
        W_PARAM = 48775;
      end
      1600: begin
        W_PARAM = 48871;
      end
      1601: begin
        W_PARAM = 15907;
      end
      1602: begin
        W_PARAM = 16006;
      end
      1603: begin
        W_PARAM = 15819;
      end
      1604: begin
        W_PARAM = 15849;
      end
      1605: begin
        W_PARAM = 16180;
      end
      1606: begin
        W_PARAM = 15548;
      end
      1607: begin
        W_PARAM = 49043;
      end
      1608: begin
        W_PARAM = 16139;
      end
      1609: begin
        W_PARAM = 48794;
      end
      1610: begin
        W_PARAM = 48648;
      end
      1611: begin
        W_PARAM = 16101;
      end
      1612: begin
        W_PARAM = 15956;
      end
      1613: begin
        W_PARAM = 48658;
      end
      1614: begin
        W_PARAM = 48398;
      end
      1615: begin
        W_PARAM = 15862;
      end
      1616: begin
        W_PARAM = 16079;
      end
      1617: begin
        W_PARAM = 48915;
      end
      1618: begin
        W_PARAM = 15873;
      end
      1619: begin
        W_PARAM = 48857;
      end
      1620: begin
        W_PARAM = 15882;
      end
      1621: begin
        W_PARAM = 16149;
      end
      1622: begin
        W_PARAM = 15829;
      end
      1623: begin
        W_PARAM = 15925;
      end
      1624: begin
        W_PARAM = 15911;
      end
      1625: begin
        W_PARAM = 16141;
      end
      1626: begin
        W_PARAM = 48878;
      end
      1627: begin
        W_PARAM = 48869;
      end
      1628: begin
        W_PARAM = 15620;
      end
      1629: begin
        W_PARAM = 48981;
      end
      1630: begin
        W_PARAM = 48870;
      end
      1631: begin
        W_PARAM = 15802;
      end
      1632: begin
        W_PARAM = 48535;
      end
      1633: begin
        W_PARAM = 48865;
      end
      1634: begin
        W_PARAM = 16205;
      end
      1635: begin
        W_PARAM = 16077;
      end
      1636: begin
        W_PARAM = 16236;
      end
      1637: begin
        W_PARAM = 48773;
      end
      1638: begin
        W_PARAM = 48863;
      end
      1639: begin
        W_PARAM = 48909;
      end
      1640: begin
        W_PARAM = 48921;
      end
      1641: begin
        W_PARAM = 48663;
      end
      1642: begin
        W_PARAM = 48910;
      end
      1643: begin
        W_PARAM = 48692;
      end
      1644: begin
        W_PARAM = 15776;
      end
      1645: begin
        W_PARAM = 16217;
      end
      1646: begin
        W_PARAM = 16085;
      end
      1647: begin
        W_PARAM = 48446;
      end
      1648: begin
        W_PARAM = 16071;
      end
      1649: begin
        W_PARAM = 48723;
      end
      1650: begin
        W_PARAM = 48786;
      end
      1651: begin
        W_PARAM = 48947;
      end
      1652: begin
        W_PARAM = 48606;
      end
      1653: begin
        W_PARAM = 48438;
      end
      1654: begin
        W_PARAM = 48716;
      end
      1655: begin
        W_PARAM = 16187;
      end
      1656: begin
        W_PARAM = 48436;
      end
      1657: begin
        W_PARAM = 48251;
      end
      1658: begin
        W_PARAM = 16189;
      end
      1659: begin
        W_PARAM = 48541;
      end
      1660: begin
        W_PARAM = 48557;
      end
      1661: begin
        W_PARAM = 48732;
      end
      1662: begin
        W_PARAM = 48506;
      end
      1663: begin
        W_PARAM = 47883;
      end
      1664: begin
        W_PARAM = 48648;
      end
      1665: begin
        W_PARAM = 15987;
      end
      1666: begin
        W_PARAM = 15988;
      end
      1667: begin
        W_PARAM = 48180;
      end
      1668: begin
        W_PARAM = 15640;
      end
      1669: begin
        W_PARAM = 48117;
      end
      1670: begin
        W_PARAM = 48415;
      end
      1671: begin
        W_PARAM = 48539;
      end
      1672: begin
        W_PARAM = 48329;
      end
      1673: begin
        W_PARAM = 47140;
      end
      1674: begin
        W_PARAM = 47619;
      end
      1675: begin
        W_PARAM = 15558;
      end
      1676: begin
        W_PARAM = 15877;
      end
      1677: begin
        W_PARAM = 47377;
      end
      1678: begin
        W_PARAM = 48235;
      end
      1679: begin
        W_PARAM = 46770;
      end
      1680: begin
        W_PARAM = 0;
      end
      1681: begin
        W_PARAM = 0;
      end
      1682: begin
        W_PARAM = 0;
      end
      1683: begin
        W_PARAM = 0;
      end
      1684: begin
        W_PARAM = 0;
      end
      1685: begin
        W_PARAM = 0;
      end
      1686: begin
        W_PARAM = 0;
      end
      1687: begin
        W_PARAM = 0;
      end
      1688: begin
        W_PARAM = 0;
      end
      1689: begin
        W_PARAM = 0;
      end
      1690: begin
        W_PARAM = 46869;
      end
      1691: begin
        W_PARAM = 46541;
      end
      1692: begin
        W_PARAM = 47503;
      end
      1693: begin
        W_PARAM = 15198;
      end
      1694: begin
        W_PARAM = 46615;
      end
      1695: begin
        W_PARAM = 47337;
      end
      1696: begin
        W_PARAM = 46155;
      end
      1697: begin
        W_PARAM = 47097;
      end
      1698: begin
        W_PARAM = 47497;
      end
      1699: begin
        W_PARAM = 47920;
      end
      1700: begin
        W_PARAM = 48087;
      end
      1701: begin
        W_PARAM = 48623;
      end
      1702: begin
        W_PARAM = 48387;
      end
      1703: begin
        W_PARAM = 15489;
      end
      1704: begin
        W_PARAM = 47995;
      end
      1705: begin
        W_PARAM = 15626;
      end
      1706: begin
        W_PARAM = 48008;
      end
      1707: begin
        W_PARAM = 15888;
      end
      1708: begin
        W_PARAM = 48270;
      end
      1709: begin
        W_PARAM = 48151;
      end
      1710: begin
        W_PARAM = 48147;
      end
      1711: begin
        W_PARAM = 15656;
      end
      1712: begin
        W_PARAM = 48095;
      end
      1713: begin
        W_PARAM = 16082;
      end
      1714: begin
        W_PARAM = 48686;
      end
      1715: begin
        W_PARAM = 48864;
      end
      1716: begin
        W_PARAM = 48676;
      end
      1717: begin
        W_PARAM = 16142;
      end
      1718: begin
        W_PARAM = 48668;
      end
      1719: begin
        W_PARAM = 48526;
      end
      1720: begin
        W_PARAM = 48592;
      end
      1721: begin
        W_PARAM = 15849;
      end
      1722: begin
        W_PARAM = 15999;
      end
      1723: begin
        W_PARAM = 15960;
      end
      1724: begin
        W_PARAM = 15564;
      end
      1725: begin
        W_PARAM = 48833;
      end
      1726: begin
        W_PARAM = 15898;
      end
      1727: begin
        W_PARAM = 16013;
      end
      1728: begin
        W_PARAM = 48811;
      end
      1729: begin
        W_PARAM = 48729;
      end
      1730: begin
        W_PARAM = 48524;
      end
      1731: begin
        W_PARAM = 15753;
      end
      1732: begin
        W_PARAM = 48556;
      end
      1733: begin
        W_PARAM = 15883;
      end
      1734: begin
        W_PARAM = 16119;
      end
      1735: begin
        W_PARAM = 15824;
      end
      1736: begin
        W_PARAM = 48730;
      end
      1737: begin
        W_PARAM = 16157;
      end
      1738: begin
        W_PARAM = 48786;
      end
      1739: begin
        W_PARAM = 48960;
      end
      1740: begin
        W_PARAM = 15886;
      end
      1741: begin
        W_PARAM = 48534;
      end
      1742: begin
        W_PARAM = 15926;
      end
      1743: begin
        W_PARAM = 16044;
      end
      1744: begin
        W_PARAM = 48513;
      end
      1745: begin
        W_PARAM = 15631;
      end
      1746: begin
        W_PARAM = 48927;
      end
      1747: begin
        W_PARAM = 16229;
      end
      1748: begin
        W_PARAM = 48803;
      end
      1749: begin
        W_PARAM = 48897;
      end
      1750: begin
        W_PARAM = 15901;
      end
      1751: begin
        W_PARAM = 48870;
      end
      1752: begin
        W_PARAM = 16032;
      end
      1753: begin
        W_PARAM = 48498;
      end
      1754: begin
        W_PARAM = 48238;
      end
      1755: begin
        W_PARAM = 48594;
      end
      1756: begin
        W_PARAM = 15767;
      end
      1757: begin
        W_PARAM = 16109;
      end
      1758: begin
        W_PARAM = 15824;
      end
      1759: begin
        W_PARAM = 48885;
      end
      1760: begin
        W_PARAM = 48258;
      end
      1761: begin
        W_PARAM = 48865;
      end
      1762: begin
        W_PARAM = 15607;
      end
      1763: begin
        W_PARAM = 16036;
      end
      1764: begin
        W_PARAM = 48752;
      end
      1765: begin
        W_PARAM = 48775;
      end
      1766: begin
        W_PARAM = 48585;
      end
      1767: begin
        W_PARAM = 16200;
      end
      1768: begin
        W_PARAM = 48580;
      end
      1769: begin
        W_PARAM = 15470;
      end
      1770: begin
        W_PARAM = 49000;
      end
      1771: begin
        W_PARAM = 48985;
      end
      1772: begin
        W_PARAM = 16116;
      end
      1773: begin
        W_PARAM = 16119;
      end
      1774: begin
        W_PARAM = 16054;
      end
      1775: begin
        W_PARAM = 48650;
      end
      1776: begin
        W_PARAM = 48788;
      end
      1777: begin
        W_PARAM = 16055;
      end
      1778: begin
        W_PARAM = 15915;
      end
      1779: begin
        W_PARAM = 16044;
      end
      1780: begin
        W_PARAM = 48746;
      end
      1781: begin
        W_PARAM = 48722;
      end
      1782: begin
        W_PARAM = 16153;
      end
      1783: begin
        W_PARAM = 16142;
      end
      1784: begin
        W_PARAM = 48834;
      end
      1785: begin
        W_PARAM = 15685;
      end
      1786: begin
        W_PARAM = 48930;
      end
      1787: begin
        W_PARAM = 16136;
      end
      1788: begin
        W_PARAM = 48523;
      end
      1789: begin
        W_PARAM = 48736;
      end
      1790: begin
        W_PARAM = 48280;
      end
      1791: begin
        W_PARAM = 15955;
      end
      1792: begin
        W_PARAM = 48733;
      end
      1793: begin
        W_PARAM = 15965;
      end
      1794: begin
        W_PARAM = 48902;
      end
      1795: begin
        W_PARAM = 48752;
      end
      1796: begin
        W_PARAM = 48859;
      end
      1797: begin
        W_PARAM = 16198;
      end
      1798: begin
        W_PARAM = 48738;
      end
      1799: begin
        W_PARAM = 16100;
      end
      1800: begin
        W_PARAM = 48920;
      end
      1801: begin
        W_PARAM = 48785;
      end
      1802: begin
        W_PARAM = 16007;
      end
      1803: begin
        W_PARAM = 48688;
      end
      1804: begin
        W_PARAM = 48750;
      end
      1805: begin
        W_PARAM = 15415;
      end
      1806: begin
        W_PARAM = 48735;
      end
      1807: begin
        W_PARAM = 16121;
      end
      1808: begin
        W_PARAM = 16159;
      end
      1809: begin
        W_PARAM = 15855;
      end
      1810: begin
        W_PARAM = 16179;
      end
      1811: begin
        W_PARAM = 48867;
      end
      1812: begin
        W_PARAM = 15183;
      end
      1813: begin
        W_PARAM = 16157;
      end
      1814: begin
        W_PARAM = 48917;
      end
      1815: begin
        W_PARAM = 48631;
      end
      1816: begin
        W_PARAM = 48954;
      end
      1817: begin
        W_PARAM = 48419;
      end
      1818: begin
        W_PARAM = 48332;
      end
      1819: begin
        W_PARAM = 16160;
      end
      1820: begin
        W_PARAM = 16063;
      end
      1821: begin
        W_PARAM = 48792;
      end
      1822: begin
        W_PARAM = 48623;
      end
      1823: begin
        W_PARAM = 15341;
      end
      1824: begin
        W_PARAM = 48922;
      end
      1825: begin
        W_PARAM = 16062;
      end
      1826: begin
        W_PARAM = 48899;
      end
      1827: begin
        W_PARAM = 15728;
      end
      1828: begin
        W_PARAM = 15812;
      end
      1829: begin
        W_PARAM = 16160;
      end
      1830: begin
        W_PARAM = 48616;
      end
      1831: begin
        W_PARAM = 48868;
      end
      1832: begin
        W_PARAM = 15963;
      end
      1833: begin
        W_PARAM = 15960;
      end
      1834: begin
        W_PARAM = 48964;
      end
      1835: begin
        W_PARAM = 48538;
      end
      1836: begin
        W_PARAM = 48287;
      end
      1837: begin
        W_PARAM = 16013;
      end
      1838: begin
        W_PARAM = 16101;
      end
      1839: begin
        W_PARAM = 16011;
      end
      1840: begin
        W_PARAM = 16040;
      end
      1841: begin
        W_PARAM = 48793;
      end
      1842: begin
        W_PARAM = 15945;
      end
      1843: begin
        W_PARAM = 16055;
      end
      1844: begin
        W_PARAM = 48937;
      end
      1845: begin
        W_PARAM = 48732;
      end
      1846: begin
        W_PARAM = 48827;
      end
      1847: begin
        W_PARAM = 15905;
      end
      1848: begin
        W_PARAM = 48594;
      end
      1849: begin
        W_PARAM = 16154;
      end
      1850: begin
        W_PARAM = 15710;
      end
      1851: begin
        W_PARAM = 48966;
      end
      1852: begin
        W_PARAM = 48590;
      end
      1853: begin
        W_PARAM = 48662;
      end
      1854: begin
        W_PARAM = 48729;
      end
      1855: begin
        W_PARAM = 15425;
      end
      1856: begin
        W_PARAM = 48639;
      end
      1857: begin
        W_PARAM = 16067;
      end
      1858: begin
        W_PARAM = 16034;
      end
      1859: begin
        W_PARAM = 16152;
      end
      1860: begin
        W_PARAM = 16126;
      end
      1861: begin
        W_PARAM = 15643;
      end
      1862: begin
        W_PARAM = 48354;
      end
      1863: begin
        W_PARAM = 16184;
      end
      1864: begin
        W_PARAM = 48968;
      end
      1865: begin
        W_PARAM = 15470;
      end
      1866: begin
        W_PARAM = 49007;
      end
      1867: begin
        W_PARAM = 16031;
      end
      1868: begin
        W_PARAM = 48830;
      end
      1869: begin
        W_PARAM = 16137;
      end
      1870: begin
        W_PARAM = 48733;
      end
      1871: begin
        W_PARAM = 48898;
      end
      1872: begin
        W_PARAM = 48379;
      end
      1873: begin
        W_PARAM = 48878;
      end
      1874: begin
        W_PARAM = 48673;
      end
      1875: begin
        W_PARAM = 16147;
      end
      1876: begin
        W_PARAM = 48817;
      end
      1877: begin
        W_PARAM = 15801;
      end
      1878: begin
        W_PARAM = 16221;
      end
      1879: begin
        W_PARAM = 15943;
      end
      1880: begin
        W_PARAM = 16030;
      end
      1881: begin
        W_PARAM = 48523;
      end
      1882: begin
        W_PARAM = 48818;
      end
      1883: begin
        W_PARAM = 16006;
      end
      1884: begin
        W_PARAM = 48897;
      end
      1885: begin
        W_PARAM = 16020;
      end
      1886: begin
        W_PARAM = 48664;
      end
      1887: begin
        W_PARAM = 48532;
      end
      1888: begin
        W_PARAM = 15387;
      end
      1889: begin
        W_PARAM = 16012;
      end
      1890: begin
        W_PARAM = 16165;
      end
      1891: begin
        W_PARAM = 48661;
      end
      1892: begin
        W_PARAM = 48740;
      end
      1893: begin
        W_PARAM = 15988;
      end
      1894: begin
        W_PARAM = 48797;
      end
      1895: begin
        W_PARAM = 48689;
      end
      1896: begin
        W_PARAM = 15492;
      end
      1897: begin
        W_PARAM = 15918;
      end
      1898: begin
        W_PARAM = 48663;
      end
      1899: begin
        W_PARAM = 48539;
      end
      1900: begin
        W_PARAM = 16238;
      end
      1901: begin
        W_PARAM = 48086;
      end
      1902: begin
        W_PARAM = 48798;
      end
      1903: begin
        W_PARAM = 48391;
      end
      1904: begin
        W_PARAM = 48460;
      end
      1905: begin
        W_PARAM = 16046;
      end
      1906: begin
        W_PARAM = 48520;
      end
      1907: begin
        W_PARAM = 48775;
      end
      1908: begin
        W_PARAM = 48649;
      end
      1909: begin
        W_PARAM = 48849;
      end
      1910: begin
        W_PARAM = 15698;
      end
      1911: begin
        W_PARAM = 16024;
      end
      1912: begin
        W_PARAM = 48970;
      end
      1913: begin
        W_PARAM = 48518;
      end
      1914: begin
        W_PARAM = 16189;
      end
      1915: begin
        W_PARAM = 15415;
      end
      1916: begin
        W_PARAM = 16100;
      end
      1917: begin
        W_PARAM = 48973;
      end
      1918: begin
        W_PARAM = 16136;
      end
      1919: begin
        W_PARAM = 48851;
      end
      1920: begin
        W_PARAM = 49009;
      end
      1921: begin
        W_PARAM = 15872;
      end
      1922: begin
        W_PARAM = 48888;
      end
      1923: begin
        W_PARAM = 15791;
      end
      1924: begin
        W_PARAM = 15627;
      end
      1925: begin
        W_PARAM = 16299;
      end
      1926: begin
        W_PARAM = 16111;
      end
      1927: begin
        W_PARAM = 48697;
      end
      1928: begin
        W_PARAM = 48473;
      end
      1929: begin
        W_PARAM = 48838;
      end
      1930: begin
        W_PARAM = 48954;
      end
      1931: begin
        W_PARAM = 48840;
      end
      1932: begin
        W_PARAM = 48481;
      end
      1933: begin
        W_PARAM = 48625;
      end
      1934: begin
        W_PARAM = 48521;
      end
      1935: begin
        W_PARAM = 16165;
      end
      1936: begin
        W_PARAM = 15741;
      end
      1937: begin
        W_PARAM = 48563;
      end
      1938: begin
        W_PARAM = 16221;
      end
      1939: begin
        W_PARAM = 48642;
      end
      1940: begin
        W_PARAM = 48831;
      end
      1941: begin
        W_PARAM = 48619;
      end
      1942: begin
        W_PARAM = 48299;
      end
      1943: begin
        W_PARAM = 48109;
      end
      1944: begin
        W_PARAM = 16019;
      end
      1945: begin
        W_PARAM = 16008;
      end
      1946: begin
        W_PARAM = 48658;
      end
      1947: begin
        W_PARAM = 48279;
      end
      1948: begin
        W_PARAM = 15929;
      end
      1949: begin
        W_PARAM = 48481;
      end
      1950: begin
        W_PARAM = 48583;
      end
      1951: begin
        W_PARAM = 47043;
      end
      1952: begin
        W_PARAM = 47439;
      end
      1953: begin
        W_PARAM = 47311;
      end
      1954: begin
        W_PARAM = 48087;
      end
      1955: begin
        W_PARAM = 15895;
      end
      1956: begin
        W_PARAM = 48276;
      end
      1957: begin
        W_PARAM = 47576;
      end
      1958: begin
        W_PARAM = 48328;
      end
      1959: begin
        W_PARAM = 47457;
      end
      1960: begin
        W_PARAM = 0;
      end
      1961: begin
        W_PARAM = 0;
      end
      1962: begin
        W_PARAM = 0;
      end
      1963: begin
        W_PARAM = 0;
      end
      1964: begin
        W_PARAM = 0;
      end
      1965: begin
        W_PARAM = 0;
      end
      1966: begin
        W_PARAM = 0;
      end
      1967: begin
        W_PARAM = 0;
      end
      1968: begin
        W_PARAM = 0;
      end
      1969: begin
        W_PARAM = 0;
      end
      1970: begin
        W_PARAM = 47662;
      end
      1971: begin
        W_PARAM = 48257;
      end
      1972: begin
        W_PARAM = 48121;
      end
      1973: begin
        W_PARAM = 15805;
      end
      1974: begin
        W_PARAM = 48006;
      end
      1975: begin
        W_PARAM = 47964;
      end
      1976: begin
        W_PARAM = 46731;
      end
      1977: begin
        W_PARAM = 15602;
      end
      1978: begin
        W_PARAM = 48272;
      end
      1979: begin
        W_PARAM = 48533;
      end
      1980: begin
        W_PARAM = 47326;
      end
      1981: begin
        W_PARAM = 48772;
      end
      1982: begin
        W_PARAM = 15932;
      end
      1983: begin
        W_PARAM = 48577;
      end
      1984: begin
        W_PARAM = 48091;
      end
      1985: begin
        W_PARAM = 48390;
      end
      1986: begin
        W_PARAM = 48280;
      end
      1987: begin
        W_PARAM = 16017;
      end
      1988: begin
        W_PARAM = 48298;
      end
      1989: begin
        W_PARAM = 48403;
      end
      1990: begin
        W_PARAM = 48177;
      end
      1991: begin
        W_PARAM = 48513;
      end
      1992: begin
        W_PARAM = 15944;
      end
      1993: begin
        W_PARAM = 15731;
      end
      1994: begin
        W_PARAM = 48464;
      end
      1995: begin
        W_PARAM = 48858;
      end
      1996: begin
        W_PARAM = 48700;
      end
      1997: begin
        W_PARAM = 16222;
      end
      1998: begin
        W_PARAM = 48667;
      end
      1999: begin
        W_PARAM = 48754;
      end
      2000: begin
        W_PARAM = 48723;
      end
      2001: begin
        W_PARAM = 15840;
      end
      2002: begin
        W_PARAM = 16211;
      end
      2003: begin
        W_PARAM = 16101;
      end
      2004: begin
        W_PARAM = 16009;
      end
      2005: begin
        W_PARAM = 49045;
      end
      2006: begin
        W_PARAM = 15913;
      end
      2007: begin
        W_PARAM = 16026;
      end
      2008: begin
        W_PARAM = 48638;
      end
      2009: begin
        W_PARAM = 48927;
      end
      2010: begin
        W_PARAM = 15578;
      end
      2011: begin
        W_PARAM = 48848;
      end
      2012: begin
        W_PARAM = 15937;
      end
      2013: begin
        W_PARAM = 16238;
      end
      2014: begin
        W_PARAM = 16236;
      end
      2015: begin
        W_PARAM = 48738;
      end
      2016: begin
        W_PARAM = 15635;
      end
      2017: begin
        W_PARAM = 48792;
      end
      2018: begin
        W_PARAM = 48474;
      end
      2019: begin
        W_PARAM = 49040;
      end
      2020: begin
        W_PARAM = 16073;
      end
      2021: begin
        W_PARAM = 48911;
      end
      2022: begin
        W_PARAM = 16190;
      end
      2023: begin
        W_PARAM = 16066;
      end
      2024: begin
        W_PARAM = 15897;
      end
      2025: begin
        W_PARAM = 48611;
      end
      2026: begin
        W_PARAM = 48978;
      end
      2027: begin
        W_PARAM = 16060;
      end
      2028: begin
        W_PARAM = 48796;
      end
      2029: begin
        W_PARAM = 48754;
      end
      2030: begin
        W_PARAM = 15755;
      end
      2031: begin
        W_PARAM = 48798;
      end
      2032: begin
        W_PARAM = 48835;
      end
      2033: begin
        W_PARAM = 15772;
      end
      2034: begin
        W_PARAM = 16035;
      end
      2035: begin
        W_PARAM = 15970;
      end
      2036: begin
        W_PARAM = 16033;
      end
      2037: begin
        W_PARAM = 16014;
      end
      2038: begin
        W_PARAM = 48737;
      end
      2039: begin
        W_PARAM = 48828;
      end
      2040: begin
        W_PARAM = 48859;
      end
      2041: begin
        W_PARAM = 49013;
      end
      2042: begin
        W_PARAM = 16132;
      end
      2043: begin
        W_PARAM = 16002;
      end
      2044: begin
        W_PARAM = 48419;
      end
      2045: begin
        W_PARAM = 16150;
      end
      2046: begin
        W_PARAM = 48773;
      end
      2047: begin
        W_PARAM = 48541;
      end
      2048: begin
        W_PARAM = 16137;
      end
      2049: begin
        W_PARAM = 48645;
      end
      2050: begin
        W_PARAM = 15924;
      end
      2051: begin
        W_PARAM = 48767;
      end
      2052: begin
        W_PARAM = 48484;
      end
      2053: begin
        W_PARAM = 15762;
      end
      2054: begin
        W_PARAM = 15904;
      end
      2055: begin
        W_PARAM = 48207;
      end
      2056: begin
        W_PARAM = 48546;
      end
      2057: begin
        W_PARAM = 16069;
      end
      2058: begin
        W_PARAM = 48706;
      end
      2059: begin
        W_PARAM = 48718;
      end
      2060: begin
        W_PARAM = 48491;
      end
      2061: begin
        W_PARAM = 16011;
      end
      2062: begin
        W_PARAM = 48804;
      end
      2063: begin
        W_PARAM = 48269;
      end
      2064: begin
        W_PARAM = 48897;
      end
      2065: begin
        W_PARAM = 16073;
      end
      2066: begin
        W_PARAM = 48806;
      end
      2067: begin
        W_PARAM = 16123;
      end
      2068: begin
        W_PARAM = 15945;
      end
      2069: begin
        W_PARAM = 48643;
      end
      2070: begin
        W_PARAM = 16098;
      end
      2071: begin
        W_PARAM = 48887;
      end
      2072: begin
        W_PARAM = 15954;
      end
      2073: begin
        W_PARAM = 48648;
      end
      2074: begin
        W_PARAM = 15831;
      end
      2075: begin
        W_PARAM = 15742;
      end
      2076: begin
        W_PARAM = 48547;
      end
      2077: begin
        W_PARAM = 16000;
      end
      2078: begin
        W_PARAM = 48825;
      end
      2079: begin
        W_PARAM = 48165;
      end
      2080: begin
        W_PARAM = 48719;
      end
      2081: begin
        W_PARAM = 16010;
      end
      2082: begin
        W_PARAM = 48777;
      end
      2083: begin
        W_PARAM = 16014;
      end
      2084: begin
        W_PARAM = 48961;
      end
      2085: begin
        W_PARAM = 15991;
      end
      2086: begin
        W_PARAM = 48655;
      end
      2087: begin
        W_PARAM = 16031;
      end
      2088: begin
        W_PARAM = 48784;
      end
      2089: begin
        W_PARAM = 16140;
      end
      2090: begin
        W_PARAM = 16003;
      end
      2091: begin
        W_PARAM = 48896;
      end
      2092: begin
        W_PARAM = 16147;
      end
      2093: begin
        W_PARAM = 48801;
      end
      2094: begin
        W_PARAM = 48696;
      end
      2095: begin
        W_PARAM = 48919;
      end
      2096: begin
        W_PARAM = 48896;
      end
      2097: begin
        W_PARAM = 16105;
      end
      2098: begin
        W_PARAM = 48144;
      end
      2099: begin
        W_PARAM = 16207;
      end
      2100: begin
        W_PARAM = 15356;
      end
      2101: begin
        W_PARAM = 48540;
      end
      2102: begin
        W_PARAM = 15734;
      end
      2103: begin
        W_PARAM = 16155;
      end
      2104: begin
        W_PARAM = 48919;
      end
      2105: begin
        W_PARAM = 16104;
      end
      2106: begin
        W_PARAM = 15875;
      end
      2107: begin
        W_PARAM = 48768;
      end
      2108: begin
        W_PARAM = 48939;
      end
      2109: begin
        W_PARAM = 16039;
      end
      2110: begin
        W_PARAM = 48756;
      end
      2111: begin
        W_PARAM = 48933;
      end
      2112: begin
        W_PARAM = 48731;
      end
      2113: begin
        W_PARAM = 16015;
      end
      2114: begin
        W_PARAM = 48775;
      end
      2115: begin
        W_PARAM = 48848;
      end
      2116: begin
        W_PARAM = 48593;
      end
      2117: begin
        W_PARAM = 16027;
      end
      2118: begin
        W_PARAM = 16140;
      end
      2119: begin
        W_PARAM = 16190;
      end
      2120: begin
        W_PARAM = 48670;
      end
      2121: begin
        W_PARAM = 48564;
      end
      2122: begin
        W_PARAM = 15346;
      end
      2123: begin
        W_PARAM = 48515;
      end
      2124: begin
        W_PARAM = 48890;
      end
      2125: begin
        W_PARAM = 16032;
      end
      2126: begin
        W_PARAM = 48924;
      end
      2127: begin
        W_PARAM = 16092;
      end
      2128: begin
        W_PARAM = 15739;
      end
      2129: begin
        W_PARAM = 16152;
      end
      2130: begin
        W_PARAM = 16127;
      end
      2131: begin
        W_PARAM = 48773;
      end
      2132: begin
        W_PARAM = 48906;
      end
      2133: begin
        W_PARAM = 16073;
      end
      2134: begin
        W_PARAM = 15888;
      end
      2135: begin
        W_PARAM = 15064;
      end
      2136: begin
        W_PARAM = 48804;
      end
      2137: begin
        W_PARAM = 16045;
      end
      2138: begin
        W_PARAM = 48905;
      end
      2139: begin
        W_PARAM = 16018;
      end
      2140: begin
        W_PARAM = 16110;
      end
      2141: begin
        W_PARAM = 48863;
      end
      2142: begin
        W_PARAM = 15872;
      end
      2143: begin
        W_PARAM = 48896;
      end
      2144: begin
        W_PARAM = 48852;
      end
      2145: begin
        W_PARAM = 15982;
      end
      2146: begin
        W_PARAM = 48840;
      end
      2147: begin
        W_PARAM = 16128;
      end
      2148: begin
        W_PARAM = 16035;
      end
      2149: begin
        W_PARAM = 15826;
      end
      2150: begin
        W_PARAM = 15963;
      end
      2151: begin
        W_PARAM = 48424;
      end
      2152: begin
        W_PARAM = 48779;
      end
      2153: begin
        W_PARAM = 16062;
      end
      2154: begin
        W_PARAM = 15872;
      end
      2155: begin
        W_PARAM = 15439;
      end
      2156: begin
        W_PARAM = 48725;
      end
      2157: begin
        W_PARAM = 15887;
      end
      2158: begin
        W_PARAM = 48815;
      end
      2159: begin
        W_PARAM = 14701;
      end
      2160: begin
        W_PARAM = 48486;
      end
      2161: begin
        W_PARAM = 15909;
      end
      2162: begin
        W_PARAM = 48892;
      end
      2163: begin
        W_PARAM = 15734;
      end
      2164: begin
        W_PARAM = 15790;
      end
      2165: begin
        W_PARAM = 48505;
      end
      2166: begin
        W_PARAM = 48942;
      end
      2167: begin
        W_PARAM = 16182;
      end
      2168: begin
        W_PARAM = 48658;
      end
      2169: begin
        W_PARAM = 16085;
      end
      2170: begin
        W_PARAM = 48747;
      end
      2171: begin
        W_PARAM = 48538;
      end
      2172: begin
        W_PARAM = 48141;
      end
      2173: begin
        W_PARAM = 48912;
      end
      2174: begin
        W_PARAM = 15720;
      end
      2175: begin
        W_PARAM = 15980;
      end
      2176: begin
        W_PARAM = 48706;
      end
      2177: begin
        W_PARAM = 16078;
      end
      2178: begin
        W_PARAM = 16106;
      end
      2179: begin
        W_PARAM = 48556;
      end
      2180: begin
        W_PARAM = 48771;
      end
      2181: begin
        W_PARAM = 48766;
      end
      2182: begin
        W_PARAM = 16188;
      end
      2183: begin
        W_PARAM = 48910;
      end
      2184: begin
        W_PARAM = 16043;
      end
      2185: begin
        W_PARAM = 16140;
      end
      2186: begin
        W_PARAM = 48909;
      end
      2187: begin
        W_PARAM = 15859;
      end
      2188: begin
        W_PARAM = 15934;
      end
      2189: begin
        W_PARAM = 48799;
      end
      2190: begin
        W_PARAM = 16108;
      end
      2191: begin
        W_PARAM = 48777;
      end
      2192: begin
        W_PARAM = 49071;
      end
      2193: begin
        W_PARAM = 48759;
      end
      2194: begin
        W_PARAM = 16161;
      end
      2195: begin
        W_PARAM = 16070;
      end
      2196: begin
        W_PARAM = 48408;
      end
      2197: begin
        W_PARAM = 48308;
      end
      2198: begin
        W_PARAM = 16132;
      end
      2199: begin
        W_PARAM = 48489;
      end
      2200: begin
        W_PARAM = 48645;
      end
      2201: begin
        W_PARAM = 49007;
      end
      2202: begin
        W_PARAM = 49010;
      end
      2203: begin
        W_PARAM = 48645;
      end
      2204: begin
        W_PARAM = 16042;
      end
      2205: begin
        W_PARAM = 16209;
      end
      2206: begin
        W_PARAM = 16187;
      end
      2207: begin
        W_PARAM = 15670;
      end
      2208: begin
        W_PARAM = 16110;
      end
      2209: begin
        W_PARAM = 48769;
      end
      2210: begin
        W_PARAM = 48952;
      end
      2211: begin
        W_PARAM = 48922;
      end
      2212: begin
        W_PARAM = 48528;
      end
      2213: begin
        W_PARAM = 48641;
      end
      2214: begin
        W_PARAM = 15749;
      end
      2215: begin
        W_PARAM = 16337;
      end
      2216: begin
        W_PARAM = 48759;
      end
      2217: begin
        W_PARAM = 48601;
      end
      2218: begin
        W_PARAM = 16025;
      end
      2219: begin
        W_PARAM = 48644;
      end
      2220: begin
        W_PARAM = 48867;
      end
      2221: begin
        W_PARAM = 48334;
      end
      2222: begin
        W_PARAM = 48370;
      end
      2223: begin
        W_PARAM = 48035;
      end
      2224: begin
        W_PARAM = 16081;
      end
      2225: begin
        W_PARAM = 15881;
      end
      2226: begin
        W_PARAM = 48665;
      end
      2227: begin
        W_PARAM = 48198;
      end
      2228: begin
        W_PARAM = 15967;
      end
      2229: begin
        W_PARAM = 48576;
      end
      2230: begin
        W_PARAM = 48306;
      end
      2231: begin
        W_PARAM = 48113;
      end
      2232: begin
        W_PARAM = 47965;
      end
      2233: begin
        W_PARAM = 47492;
      end
      2234: begin
        W_PARAM = 48215;
      end
      2235: begin
        W_PARAM = 15762;
      end
      2236: begin
        W_PARAM = 48438;
      end
      2237: begin
        W_PARAM = 47409;
      end
      2238: begin
        W_PARAM = 15527;
      end
      2239: begin
        W_PARAM = 47802;
      end
      2240: begin
        W_PARAM = 15773;
      end
      2241: begin
        W_PARAM = 46184;
      end
      2242: begin
        W_PARAM = 47619;
      end
      2243: begin
        W_PARAM = 46227;
      end
      2244: begin
        W_PARAM = 47925;
      end
      2245: begin
        W_PARAM = 46511;
      end
      2246: begin
        W_PARAM = 46597;
      end
      2247: begin
        W_PARAM = 48481;
      end
      2248: begin
        W_PARAM = 47012;
      end
      2249: begin
        W_PARAM = 48280;
      end
      2250: begin
        W_PARAM = 47560;
      end
      2251: begin
        W_PARAM = 48213;
      end
      2252: begin
        W_PARAM = 15312;
      end
      2253: begin
        W_PARAM = 48455;
      end
      2254: begin
        W_PARAM = 48455;
      end
      2255: begin
        W_PARAM = 47746;
      end
      2256: begin
        W_PARAM = 47283;
      end
      2257: begin
        W_PARAM = 15965;
      end
      2258: begin
        W_PARAM = 48258;
      end
      2259: begin
        W_PARAM = 48578;
      end
      2260: begin
        W_PARAM = 15524;
      end
      2261: begin
        W_PARAM = 48696;
      end
      2262: begin
        W_PARAM = 15759;
      end
      2263: begin
        W_PARAM = 48542;
      end
      2264: begin
        W_PARAM = 15900;
      end
      2265: begin
        W_PARAM = 48458;
      end
      2266: begin
        W_PARAM = 48248;
      end
      2267: begin
        W_PARAM = 16009;
      end
      2268: begin
        W_PARAM = 48393;
      end
      2269: begin
        W_PARAM = 48671;
      end
      2270: begin
        W_PARAM = 15801;
      end
      2271: begin
        W_PARAM = 48173;
      end
      2272: begin
        W_PARAM = 15136;
      end
      2273: begin
        W_PARAM = 15772;
      end
      2274: begin
        W_PARAM = 15891;
      end
      2275: begin
        W_PARAM = 48878;
      end
      2276: begin
        W_PARAM = 48664;
      end
      2277: begin
        W_PARAM = 16224;
      end
      2278: begin
        W_PARAM = 15850;
      end
      2279: begin
        W_PARAM = 48942;
      end
      2280: begin
        W_PARAM = 48741;
      end
      2281: begin
        W_PARAM = 15396;
      end
      2282: begin
        W_PARAM = 16184;
      end
      2283: begin
        W_PARAM = 16075;
      end
      2284: begin
        W_PARAM = 15957;
      end
      2285: begin
        W_PARAM = 49097;
      end
      2286: begin
        W_PARAM = 15955;
      end
      2287: begin
        W_PARAM = 16145;
      end
      2288: begin
        W_PARAM = 16029;
      end
      2289: begin
        W_PARAM = 48927;
      end
      2290: begin
        W_PARAM = 48646;
      end
      2291: begin
        W_PARAM = 48727;
      end
      2292: begin
        W_PARAM = 48706;
      end
      2293: begin
        W_PARAM = 48186;
      end
      2294: begin
        W_PARAM = 16194;
      end
      2295: begin
        W_PARAM = 48831;
      end
      2296: begin
        W_PARAM = 48634;
      end
      2297: begin
        W_PARAM = 16024;
      end
      2298: begin
        W_PARAM = 16017;
      end
      2299: begin
        W_PARAM = 48793;
      end
      2300: begin
        W_PARAM = 48650;
      end
      2301: begin
        W_PARAM = 48908;
      end
      2302: begin
        W_PARAM = 48173;
      end
      2303: begin
        W_PARAM = 48632;
      end
      2304: begin
        W_PARAM = 15840;
      end
      2305: begin
        W_PARAM = 15629;
      end
      2306: begin
        W_PARAM = 48847;
      end
      2307: begin
        W_PARAM = 16024;
      end
      2308: begin
        W_PARAM = 16129;
      end
      2309: begin
        W_PARAM = 16009;
      end
      2310: begin
        W_PARAM = 48424;
      end
      2311: begin
        W_PARAM = 15877;
      end
      2312: begin
        W_PARAM = 15859;
      end
      2313: begin
        W_PARAM = 48411;
      end
      2314: begin
        W_PARAM = 15998;
      end
      2315: begin
        W_PARAM = 48897;
      end
      2316: begin
        W_PARAM = 48823;
      end
      2317: begin
        W_PARAM = 16257;
      end
      2318: begin
        W_PARAM = 16029;
      end
      2319: begin
        W_PARAM = 48992;
      end
      2320: begin
        W_PARAM = 15978;
      end
      2321: begin
        W_PARAM = 48957;
      end
      2322: begin
        W_PARAM = 15903;
      end
      2323: begin
        W_PARAM = 48736;
      end
      2324: begin
        W_PARAM = 48820;
      end
      2325: begin
        W_PARAM = 15962;
      end
      2326: begin
        W_PARAM = 48896;
      end
      2327: begin
        W_PARAM = 16173;
      end
      2328: begin
        W_PARAM = 48766;
      end
      2329: begin
        W_PARAM = 16202;
      end
      2330: begin
        W_PARAM = 16168;
      end
      2331: begin
        W_PARAM = 48976;
      end
      2332: begin
        W_PARAM = 48684;
      end
      2333: begin
        W_PARAM = 48843;
      end
      2334: begin
        W_PARAM = 16036;
      end
      2335: begin
        W_PARAM = 15858;
      end
      2336: begin
        W_PARAM = 15612;
      end
      2337: begin
        W_PARAM = 16000;
      end
      2338: begin
        W_PARAM = 15980;
      end
      2339: begin
        W_PARAM = 48744;
      end
      2340: begin
        W_PARAM = 48823;
      end
      2341: begin
        W_PARAM = 48575;
      end
      2342: begin
        W_PARAM = 16087;
      end
      2343: begin
        W_PARAM = 15934;
      end
      2344: begin
        W_PARAM = 48809;
      end
      2345: begin
        W_PARAM = 15916;
      end
      2346: begin
        W_PARAM = 48571;
      end
      2347: begin
        W_PARAM = 15595;
      end
      2348: begin
        W_PARAM = 15993;
      end
      2349: begin
        W_PARAM = 48690;
      end
      2350: begin
        W_PARAM = 48706;
      end
      2351: begin
        W_PARAM = 48909;
      end
      2352: begin
        W_PARAM = 15728;
      end
      2353: begin
        W_PARAM = 15622;
      end
      2354: begin
        W_PARAM = 16024;
      end
      2355: begin
        W_PARAM = 15709;
      end
      2356: begin
        W_PARAM = 48783;
      end
      2357: begin
        W_PARAM = 16168;
      end
      2358: begin
        W_PARAM = 47746;
      end
      2359: begin
        W_PARAM = 48538;
      end
      2360: begin
        W_PARAM = 16130;
      end
      2361: begin
        W_PARAM = 15679;
      end
      2362: begin
        W_PARAM = 48647;
      end
      2363: begin
        W_PARAM = 15887;
      end
      2364: begin
        W_PARAM = 48812;
      end
      2365: begin
        W_PARAM = 48653;
      end
      2366: begin
        W_PARAM = 48820;
      end
      2367: begin
        W_PARAM = 16134;
      end
      2368: begin
        W_PARAM = 16086;
      end
      2369: begin
        W_PARAM = 48942;
      end
      2370: begin
        W_PARAM = 48748;
      end
      2371: begin
        W_PARAM = 15714;
      end
      2372: begin
        W_PARAM = 48527;
      end
      2373: begin
        W_PARAM = 15960;
      end
      2374: begin
        W_PARAM = 48883;
      end
      2375: begin
        W_PARAM = 15600;
      end
      2376: begin
        W_PARAM = 48581;
      end
      2377: begin
        W_PARAM = 48708;
      end
      2378: begin
        W_PARAM = 16131;
      end
      2379: begin
        W_PARAM = 16004;
      end
      2380: begin
        W_PARAM = 16144;
      end
      2381: begin
        W_PARAM = 48325;
      end
      2382: begin
        W_PARAM = 48286;
      end
      2383: begin
        W_PARAM = 15887;
      end
      2384: begin
        W_PARAM = 48919;
      end
      2385: begin
        W_PARAM = 48647;
      end
      2386: begin
        W_PARAM = 48954;
      end
      2387: begin
        W_PARAM = 16137;
      end
      2388: begin
        W_PARAM = 48810;
      end
      2389: begin
        W_PARAM = 16150;
      end
      2390: begin
        W_PARAM = 16069;
      end
      2391: begin
        W_PARAM = 15776;
      end
      2392: begin
        W_PARAM = 48309;
      end
      2393: begin
        W_PARAM = 15746;
      end
      2394: begin
        W_PARAM = 48659;
      end
      2395: begin
        W_PARAM = 48783;
      end
      2396: begin
        W_PARAM = 48994;
      end
      2397: begin
        W_PARAM = 16164;
      end
      2398: begin
        W_PARAM = 48472;
      end
      2399: begin
        W_PARAM = 15961;
      end
      2400: begin
        W_PARAM = 16275;
      end
      2401: begin
        W_PARAM = 48969;
      end
      2402: begin
        W_PARAM = 48780;
      end
      2403: begin
        W_PARAM = 15906;
      end
      2404: begin
        W_PARAM = 48978;
      end
      2405: begin
        W_PARAM = 15882;
      end
      2406: begin
        W_PARAM = 48856;
      end
      2407: begin
        W_PARAM = 16031;
      end
      2408: begin
        W_PARAM = 15993;
      end
      2409: begin
        W_PARAM = 16029;
      end
      2410: begin
        W_PARAM = 16020;
      end
      2411: begin
        W_PARAM = 16103;
      end
      2412: begin
        W_PARAM = 15964;
      end
      2413: begin
        W_PARAM = 48166;
      end
      2414: begin
        W_PARAM = 48838;
      end
      2415: begin
        W_PARAM = 48440;
      end
      2416: begin
        W_PARAM = 48594;
      end
      2417: begin
        W_PARAM = 48246;
      end
      2418: begin
        W_PARAM = 48765;
      end
      2419: begin
        W_PARAM = 48664;
      end
      2420: begin
        W_PARAM = 15898;
      end
      2421: begin
        W_PARAM = 48858;
      end
      2422: begin
        W_PARAM = 48909;
      end
      2423: begin
        W_PARAM = 16164;
      end
      2424: begin
        W_PARAM = 15749;
      end
      2425: begin
        W_PARAM = 48678;
      end
      2426: begin
        W_PARAM = 48981;
      end
      2427: begin
        W_PARAM = 16197;
      end
      2428: begin
        W_PARAM = 15658;
      end
      2429: begin
        W_PARAM = 16027;
      end
      2430: begin
        W_PARAM = 48838;
      end
      2431: begin
        W_PARAM = 15647;
      end
      2432: begin
        W_PARAM = 16136;
      end
      2433: begin
        W_PARAM = 48356;
      end
      2434: begin
        W_PARAM = 48823;
      end
      2435: begin
        W_PARAM = 15887;
      end
      2436: begin
        W_PARAM = 48890;
      end
      2437: begin
        W_PARAM = 15601;
      end
      2438: begin
        W_PARAM = 16121;
      end
      2439: begin
        W_PARAM = 15618;
      end
      2440: begin
        W_PARAM = 16132;
      end
      2441: begin
        W_PARAM = 48914;
      end
      2442: begin
        W_PARAM = 15939;
      end
      2443: begin
        W_PARAM = 15771;
      end
      2444: begin
        W_PARAM = 48738;
      end
      2445: begin
        W_PARAM = 16064;
      end
      2446: begin
        W_PARAM = 48850;
      end
      2447: begin
        W_PARAM = 16128;
      end
      2448: begin
        W_PARAM = 15644;
      end
      2449: begin
        W_PARAM = 48892;
      end
      2450: begin
        W_PARAM = 16130;
      end
      2451: begin
        W_PARAM = 48865;
      end
      2452: begin
        W_PARAM = 48897;
      end
      2453: begin
        W_PARAM = 15676;
      end
      2454: begin
        W_PARAM = 15892;
      end
      2455: begin
        W_PARAM = 48603;
      end
      2456: begin
        W_PARAM = 48663;
      end
      2457: begin
        W_PARAM = 48799;
      end
      2458: begin
        W_PARAM = 16023;
      end
      2459: begin
        W_PARAM = 16132;
      end
      2460: begin
        W_PARAM = 16108;
      end
      2461: begin
        W_PARAM = 48784;
      end
      2462: begin
        W_PARAM = 48713;
      end
      2463: begin
        W_PARAM = 16260;
      end
      2464: begin
        W_PARAM = 48993;
      end
      2465: begin
        W_PARAM = 48614;
      end
      2466: begin
        W_PARAM = 48943;
      end
      2467: begin
        W_PARAM = 16116;
      end
      2468: begin
        W_PARAM = 16030;
      end
      2469: begin
        W_PARAM = 48639;
      end
      2470: begin
        W_PARAM = 16160;
      end
      2471: begin
        W_PARAM = 49021;
      end
      2472: begin
        W_PARAM = 16121;
      end
      2473: begin
        W_PARAM = 49043;
      end
      2474: begin
        W_PARAM = 16016;
      end
      2475: begin
        W_PARAM = 16266;
      end
      2476: begin
        W_PARAM = 48965;
      end
      2477: begin
        W_PARAM = 16026;
      end
      2478: begin
        W_PARAM = 16047;
      end
      2479: begin
        W_PARAM = 48722;
      end
      2480: begin
        W_PARAM = 16056;
      end
      2481: begin
        W_PARAM = 49060;
      end
      2482: begin
        W_PARAM = 49039;
      end
      2483: begin
        W_PARAM = 49013;
      end
      2484: begin
        W_PARAM = 15999;
      end
      2485: begin
        W_PARAM = 16365;
      end
      2486: begin
        W_PARAM = 48833;
      end
      2487: begin
        W_PARAM = 48714;
      end
      2488: begin
        W_PARAM = 16296;
      end
      2489: begin
        W_PARAM = 15903;
      end
      2490: begin
        W_PARAM = 49018;
      end
      2491: begin
        W_PARAM = 48929;
      end
      2492: begin
        W_PARAM = 48831;
      end
      2493: begin
        W_PARAM = 48669;
      end
      2494: begin
        W_PARAM = 16182;
      end
      2495: begin
        W_PARAM = 16333;
      end
      2496: begin
        W_PARAM = 48876;
      end
      2497: begin
        W_PARAM = 48792;
      end
      2498: begin
        W_PARAM = 16168;
      end
      2499: begin
        W_PARAM = 48552;
      end
      2500: begin
        W_PARAM = 48860;
      end
      2501: begin
        W_PARAM = 48404;
      end
      2502: begin
        W_PARAM = 48450;
      end
      2503: begin
        W_PARAM = 48050;
      end
      2504: begin
        W_PARAM = 48693;
      end
      2505: begin
        W_PARAM = 16162;
      end
      2506: begin
        W_PARAM = 48816;
      end
      2507: begin
        W_PARAM = 48382;
      end
      2508: begin
        W_PARAM = 16139;
      end
      2509: begin
        W_PARAM = 48596;
      end
      2510: begin
        W_PARAM = 48274;
      end
      2511: begin
        W_PARAM = 48052;
      end
      2512: begin
        W_PARAM = 48080;
      end
      2513: begin
        W_PARAM = 47207;
      end
      2514: begin
        W_PARAM = 48144;
      end
      2515: begin
        W_PARAM = 15336;
      end
      2516: begin
        W_PARAM = 48415;
      end
      2517: begin
        W_PARAM = 48125;
      end
      2518: begin
        W_PARAM = 15782;
      end
      2519: begin
        W_PARAM = 47941;
      end
      2520: begin
        W_PARAM = 46553;
      end
      2521: begin
        W_PARAM = 47302;
      end
      2522: begin
        W_PARAM = 46891;
      end
      2523: begin
        W_PARAM = 47501;
      end
      2524: begin
        W_PARAM = 47744;
      end
      2525: begin
        W_PARAM = 47227;
      end
      2526: begin
        W_PARAM = 46361;
      end
      2527: begin
        W_PARAM = 15267;
      end
      2528: begin
        W_PARAM = 46783;
      end
      2529: begin
        W_PARAM = 47976;
      end
      2530: begin
        W_PARAM = 47740;
      end
      2531: begin
        W_PARAM = 47735;
      end
      2532: begin
        W_PARAM = 47935;
      end
      2533: begin
        W_PARAM = 48508;
      end
      2534: begin
        W_PARAM = 48418;
      end
      2535: begin
        W_PARAM = 47837;
      end
      2536: begin
        W_PARAM = 47823;
      end
      2537: begin
        W_PARAM = 15984;
      end
      2538: begin
        W_PARAM = 48090;
      end
      2539: begin
        W_PARAM = 48627;
      end
      2540: begin
        W_PARAM = 15673;
      end
      2541: begin
        W_PARAM = 48625;
      end
      2542: begin
        W_PARAM = 48688;
      end
      2543: begin
        W_PARAM = 15936;
      end
      2544: begin
        W_PARAM = 15891;
      end
      2545: begin
        W_PARAM = 48304;
      end
      2546: begin
        W_PARAM = 48417;
      end
      2547: begin
        W_PARAM = 16026;
      end
      2548: begin
        W_PARAM = 48610;
      end
      2549: begin
        W_PARAM = 48734;
      end
      2550: begin
        W_PARAM = 15966;
      end
      2551: begin
        W_PARAM = 48367;
      end
      2552: begin
        W_PARAM = 15869;
      end
      2553: begin
        W_PARAM = 16079;
      end
      2554: begin
        W_PARAM = 48812;
      end
      2555: begin
        W_PARAM = 48901;
      end
      2556: begin
        W_PARAM = 48724;
      end
      2557: begin
        W_PARAM = 16206;
      end
      2558: begin
        W_PARAM = 15407;
      end
      2559: begin
        W_PARAM = 48879;
      end
      2560: begin
        W_PARAM = 48466;
      end
      2561: begin
        W_PARAM = 48759;
      end
      2562: begin
        W_PARAM = 16101;
      end
      2563: begin
        W_PARAM = 16275;
      end
      2564: begin
        W_PARAM = 48966;
      end
      2565: begin
        W_PARAM = 49018;
      end
      2566: begin
        W_PARAM = 16108;
      end
      2567: begin
        W_PARAM = 16172;
      end
      2568: begin
        W_PARAM = 15693;
      end
      2569: begin
        W_PARAM = 48957;
      end
      2570: begin
        W_PARAM = 48578;
      end
      2571: begin
        W_PARAM = 48958;
      end
      2572: begin
        W_PARAM = 16255;
      end
      2573: begin
        W_PARAM = 15983;
      end
      2574: begin
        W_PARAM = 15633;
      end
      2575: begin
        W_PARAM = 48848;
      end
      2576: begin
        W_PARAM = 48910;
      end
      2577: begin
        W_PARAM = 16071;
      end
      2578: begin
        W_PARAM = 15711;
      end
      2579: begin
        W_PARAM = 15807;
      end
      2580: begin
        W_PARAM = 48713;
      end
      2581: begin
        W_PARAM = 48898;
      end
      2582: begin
        W_PARAM = 48982;
      end
      2583: begin
        W_PARAM = 16010;
      end
      2584: begin
        W_PARAM = 48566;
      end
      2585: begin
        W_PARAM = 15454;
      end
      2586: begin
        W_PARAM = 48848;
      end
      2587: begin
        W_PARAM = 16168;
      end
      2588: begin
        W_PARAM = 16099;
      end
      2589: begin
        W_PARAM = 16168;
      end
      2590: begin
        W_PARAM = 48790;
      end
      2591: begin
        W_PARAM = 16001;
      end
      2592: begin
        W_PARAM = 48681;
      end
      2593: begin
        W_PARAM = 16031;
      end
      2594: begin
        W_PARAM = 48659;
      end
      2595: begin
        W_PARAM = 48570;
      end
      2596: begin
        W_PARAM = 15735;
      end
      2597: begin
        W_PARAM = 15703;
      end
      2598: begin
        W_PARAM = 15270;
      end
      2599: begin
        W_PARAM = 15419;
      end
      2600: begin
        W_PARAM = 48801;
      end
      2601: begin
        W_PARAM = 15734;
      end
      2602: begin
        W_PARAM = 48580;
      end
      2603: begin
        W_PARAM = 16015;
      end
      2604: begin
        W_PARAM = 15416;
      end
      2605: begin
        W_PARAM = 48397;
      end
      2606: begin
        W_PARAM = 48909;
      end
      2607: begin
        W_PARAM = 15980;
      end
      2608: begin
        W_PARAM = 16058;
      end
      2609: begin
        W_PARAM = 15700;
      end
      2610: begin
        W_PARAM = 15766;
      end
      2611: begin
        W_PARAM = 48914;
      end
      2612: begin
        W_PARAM = 15966;
      end
      2613: begin
        W_PARAM = 16016;
      end
      2614: begin
        W_PARAM = 48499;
      end
      2615: begin
        W_PARAM = 48833;
      end
      2616: begin
        W_PARAM = 48779;
      end
      2617: begin
        W_PARAM = 16135;
      end
      2618: begin
        W_PARAM = 15992;
      end
      2619: begin
        W_PARAM = 48502;
      end
      2620: begin
        W_PARAM = 16154;
      end
      2621: begin
        W_PARAM = 48711;
      end
      2622: begin
        W_PARAM = 16066;
      end
      2623: begin
        W_PARAM = 48627;
      end
      2624: begin
        W_PARAM = 48898;
      end
      2625: begin
        W_PARAM = 15992;
      end
      2626: begin
        W_PARAM = 48920;
      end
      2627: begin
        W_PARAM = 48668;
      end
      2628: begin
        W_PARAM = 15716;
      end
      2629: begin
        W_PARAM = 16021;
      end
      2630: begin
        W_PARAM = 48448;
      end
      2631: begin
        W_PARAM = 48782;
      end
      2632: begin
        W_PARAM = 48875;
      end
      2633: begin
        W_PARAM = 48896;
      end
      2634: begin
        W_PARAM = 15861;
      end
      2635: begin
        W_PARAM = 16086;
      end
      2636: begin
        W_PARAM = 48432;
      end
      2637: begin
        W_PARAM = 16000;
      end
      2638: begin
        W_PARAM = 15945;
      end
      2639: begin
        W_PARAM = 16048;
      end
      2640: begin
        W_PARAM = 48603;
      end
      2641: begin
        W_PARAM = 48801;
      end
      2642: begin
        W_PARAM = 15508;
      end
      2643: begin
        W_PARAM = 48699;
      end
      2644: begin
        W_PARAM = 48712;
      end
      2645: begin
        W_PARAM = 16018;
      end
      2646: begin
        W_PARAM = 48787;
      end
      2647: begin
        W_PARAM = 16260;
      end
      2648: begin
        W_PARAM = 48871;
      end
      2649: begin
        W_PARAM = 15949;
      end
      2650: begin
        W_PARAM = 16203;
      end
      2651: begin
        W_PARAM = 15872;
      end
      2652: begin
        W_PARAM = 48779;
      end
      2653: begin
        W_PARAM = 48744;
      end
      2654: begin
        W_PARAM = 15423;
      end
      2655: begin
        W_PARAM = 48544;
      end
      2656: begin
        W_PARAM = 48973;
      end
      2657: begin
        W_PARAM = 15884;
      end
      2658: begin
        W_PARAM = 15816;
      end
      2659: begin
        W_PARAM = 15958;
      end
      2660: begin
        W_PARAM = 48518;
      end
      2661: begin
        W_PARAM = 15618;
      end
      2662: begin
        W_PARAM = 48563;
      end
      2663: begin
        W_PARAM = 16064;
      end
      2664: begin
        W_PARAM = 48959;
      end
      2665: begin
        W_PARAM = 48812;
      end
      2666: begin
        W_PARAM = 48406;
      end
      2667: begin
        W_PARAM = 16264;
      end
      2668: begin
        W_PARAM = 48828;
      end
      2669: begin
        W_PARAM = 15913;
      end
      2670: begin
        W_PARAM = 48975;
      end
      2671: begin
        W_PARAM = 16183;
      end
      2672: begin
        W_PARAM = 16066;
      end
      2673: begin
        W_PARAM = 16161;
      end
      2674: begin
        W_PARAM = 48880;
      end
      2675: begin
        W_PARAM = 48910;
      end
      2676: begin
        W_PARAM = 48851;
      end
      2677: begin
        W_PARAM = 16136;
      end
      2678: begin
        W_PARAM = 48920;
      end
      2679: begin
        W_PARAM = 16151;
      end
      2680: begin
        W_PARAM = 15962;
      end
      2681: begin
        W_PARAM = 16065;
      end
      2682: begin
        W_PARAM = 16096;
      end
      2683: begin
        W_PARAM = 16042;
      end
      2684: begin
        W_PARAM = 15954;
      end
      2685: begin
        W_PARAM = 48905;
      end
      2686: begin
        W_PARAM = 49000;
      end
      2687: begin
        W_PARAM = 15920;
      end
      2688: begin
        W_PARAM = 48462;
      end
      2689: begin
        W_PARAM = 48761;
      end
      2690: begin
        W_PARAM = 15962;
      end
      2691: begin
        W_PARAM = 48652;
      end
      2692: begin
        W_PARAM = 48815;
      end
      2693: begin
        W_PARAM = 15962;
      end
      2694: begin
        W_PARAM = 48660;
      end
      2695: begin
        W_PARAM = 48714;
      end
      2696: begin
        W_PARAM = 49049;
      end
      2697: begin
        W_PARAM = 16280;
      end
      2698: begin
        W_PARAM = 15946;
      end
      2699: begin
        W_PARAM = 15954;
      end
      2700: begin
        W_PARAM = 16010;
      end
      2701: begin
        W_PARAM = 48465;
      end
      2702: begin
        W_PARAM = 15796;
      end
      2703: begin
        W_PARAM = 48304;
      end
      2704: begin
        W_PARAM = 16017;
      end
      2705: begin
        W_PARAM = 48549;
      end
      2706: begin
        W_PARAM = 48958;
      end
      2707: begin
        W_PARAM = 16003;
      end
      2708: begin
        W_PARAM = 48702;
      end
      2709: begin
        W_PARAM = 15931;
      end
      2710: begin
        W_PARAM = 16170;
      end
      2711: begin
        W_PARAM = 48776;
      end
      2712: begin
        W_PARAM = 48603;
      end
      2713: begin
        W_PARAM = 16035;
      end
      2714: begin
        W_PARAM = 48770;
      end
      2715: begin
        W_PARAM = 48660;
      end
      2716: begin
        W_PARAM = 48948;
      end
      2717: begin
        W_PARAM = 16151;
      end
      2718: begin
        W_PARAM = 48594;
      end
      2719: begin
        W_PARAM = 14930;
      end
      2720: begin
        W_PARAM = 16089;
      end
      2721: begin
        W_PARAM = 48898;
      end
      2722: begin
        W_PARAM = 48688;
      end
      2723: begin
        W_PARAM = 16077;
      end
      2724: begin
        W_PARAM = 15984;
      end
      2725: begin
        W_PARAM = 48654;
      end
      2726: begin
        W_PARAM = 48872;
      end
      2727: begin
        W_PARAM = 48653;
      end
      2728: begin
        W_PARAM = 15794;
      end
      2729: begin
        W_PARAM = 16009;
      end
      2730: begin
        W_PARAM = 48893;
      end
      2731: begin
        W_PARAM = 48684;
      end
      2732: begin
        W_PARAM = 48836;
      end
      2733: begin
        W_PARAM = 15650;
      end
      2734: begin
        W_PARAM = 15757;
      end
      2735: begin
        W_PARAM = 16153;
      end
      2736: begin
        W_PARAM = 16005;
      end
      2737: begin
        W_PARAM = 16110;
      end
      2738: begin
        W_PARAM = 16022;
      end
      2739: begin
        W_PARAM = 48941;
      end
      2740: begin
        W_PARAM = 48967;
      end
      2741: begin
        W_PARAM = 48809;
      end
      2742: begin
        W_PARAM = 15618;
      end
      2743: begin
        W_PARAM = 16243;
      end
      2744: begin
        W_PARAM = 48491;
      end
      2745: begin
        W_PARAM = 16102;
      end
      2746: begin
        W_PARAM = 48975;
      end
      2747: begin
        W_PARAM = 16034;
      end
      2748: begin
        W_PARAM = 15885;
      end
      2749: begin
        W_PARAM = 15787;
      end
      2750: begin
        W_PARAM = 16167;
      end
      2751: begin
        W_PARAM = 48983;
      end
      2752: begin
        W_PARAM = 15756;
      end
      2753: begin
        W_PARAM = 48901;
      end
      2754: begin
        W_PARAM = 16150;
      end
      2755: begin
        W_PARAM = 16155;
      end
      2756: begin
        W_PARAM = 48842;
      end
      2757: begin
        W_PARAM = 15880;
      end
      2758: begin
        W_PARAM = 15997;
      end
      2759: begin
        W_PARAM = 48907;
      end
      2760: begin
        W_PARAM = 16280;
      end
      2761: begin
        W_PARAM = 48921;
      end
      2762: begin
        W_PARAM = 49052;
      end
      2763: begin
        W_PARAM = 49043;
      end
      2764: begin
        W_PARAM = 48898;
      end
      2765: begin
        W_PARAM = 16382;
      end
      2766: begin
        W_PARAM = 48802;
      end
      2767: begin
        W_PARAM = 15680;
      end
      2768: begin
        W_PARAM = 16174;
      end
      2769: begin
        W_PARAM = 48611;
      end
      2770: begin
        W_PARAM = 48958;
      end
      2771: begin
        W_PARAM = 48862;
      end
      2772: begin
        W_PARAM = 48776;
      end
      2773: begin
        W_PARAM = 48561;
      end
      2774: begin
        W_PARAM = 48812;
      end
      2775: begin
        W_PARAM = 16355;
      end
      2776: begin
        W_PARAM = 48977;
      end
      2777: begin
        W_PARAM = 15822;
      end
      2778: begin
        W_PARAM = 16265;
      end
      2779: begin
        W_PARAM = 48774;
      end
      2780: begin
        W_PARAM = 48826;
      end
      2781: begin
        W_PARAM = 48455;
      end
      2782: begin
        W_PARAM = 15641;
      end
      2783: begin
        W_PARAM = 48393;
      end
      2784: begin
        W_PARAM = 48665;
      end
      2785: begin
        W_PARAM = 16011;
      end
      2786: begin
        W_PARAM = 48875;
      end
      2787: begin
        W_PARAM = 15887;
      end
      2788: begin
        W_PARAM = 16195;
      end
      2789: begin
        W_PARAM = 48670;
      end
      2790: begin
        W_PARAM = 47853;
      end
      2791: begin
        W_PARAM = 48054;
      end
      2792: begin
        W_PARAM = 47875;
      end
      2793: begin
        W_PARAM = 47520;
      end
      2794: begin
        W_PARAM = 48274;
      end
      2795: begin
        W_PARAM = 15380;
      end
      2796: begin
        W_PARAM = 48201;
      end
      2797: begin
        W_PARAM = 16018;
      end
      2798: begin
        W_PARAM = 48764;
      end
      2799: begin
        W_PARAM = 48148;
      end
      2800: begin
        W_PARAM = 46596;
      end
      2801: begin
        W_PARAM = 47334;
      end
      2802: begin
        W_PARAM = 47025;
      end
      2803: begin
        W_PARAM = 47626;
      end
      2804: begin
        W_PARAM = 47765;
      end
      2805: begin
        W_PARAM = 47254;
      end
      2806: begin
        W_PARAM = 46386;
      end
      2807: begin
        W_PARAM = 15306;
      end
      2808: begin
        W_PARAM = 46833;
      end
      2809: begin
        W_PARAM = 48012;
      end
      2810: begin
        W_PARAM = 47632;
      end
      2811: begin
        W_PARAM = 47624;
      end
      2812: begin
        W_PARAM = 47803;
      end
      2813: begin
        W_PARAM = 48445;
      end
      2814: begin
        W_PARAM = 48411;
      end
      2815: begin
        W_PARAM = 47839;
      end
      2816: begin
        W_PARAM = 47701;
      end
      2817: begin
        W_PARAM = 15960;
      end
      2818: begin
        W_PARAM = 47976;
      end
      2819: begin
        W_PARAM = 48627;
      end
      2820: begin
        W_PARAM = 15947;
      end
      2821: begin
        W_PARAM = 48500;
      end
      2822: begin
        W_PARAM = 48637;
      end
      2823: begin
        W_PARAM = 15340;
      end
      2824: begin
        W_PARAM = 48323;
      end
      2825: begin
        W_PARAM = 48376;
      end
      2826: begin
        W_PARAM = 48669;
      end
      2827: begin
        W_PARAM = 16157;
      end
      2828: begin
        W_PARAM = 48532;
      end
      2829: begin
        W_PARAM = 48821;
      end
      2830: begin
        W_PARAM = 15899;
      end
      2831: begin
        W_PARAM = 48712;
      end
      2832: begin
        W_PARAM = 16098;
      end
      2833: begin
        W_PARAM = 16203;
      end
      2834: begin
        W_PARAM = 48682;
      end
      2835: begin
        W_PARAM = 48918;
      end
      2836: begin
        W_PARAM = 48760;
      end
      2837: begin
        W_PARAM = 16056;
      end
      2838: begin
        W_PARAM = 48812;
      end
      2839: begin
        W_PARAM = 48733;
      end
      2840: begin
        W_PARAM = 15774;
      end
      2841: begin
        W_PARAM = 48839;
      end
      2842: begin
        W_PARAM = 48826;
      end
      2843: begin
        W_PARAM = 16056;
      end
      2844: begin
        W_PARAM = 48828;
      end
      2845: begin
        W_PARAM = 48570;
      end
      2846: begin
        W_PARAM = 48319;
      end
      2847: begin
        W_PARAM = 16107;
      end
      2848: begin
        W_PARAM = 16191;
      end
      2849: begin
        W_PARAM = 48848;
      end
      2850: begin
        W_PARAM = 16117;
      end
      2851: begin
        W_PARAM = 48967;
      end
      2852: begin
        W_PARAM = 16252;
      end
      2853: begin
        W_PARAM = 48675;
      end
      2854: begin
        W_PARAM = 48800;
      end
      2855: begin
        W_PARAM = 48483;
      end
      2856: begin
        W_PARAM = 48863;
      end
      2857: begin
        W_PARAM = 16013;
      end
      2858: begin
        W_PARAM = 48649;
      end
      2859: begin
        W_PARAM = 15883;
      end
      2860: begin
        W_PARAM = 48200;
      end
      2861: begin
        W_PARAM = 49040;
      end
      2862: begin
        W_PARAM = 16246;
      end
      2863: begin
        W_PARAM = 15975;
      end
      2864: begin
        W_PARAM = 48897;
      end
      2865: begin
        W_PARAM = 48908;
      end
      2866: begin
        W_PARAM = 48721;
      end
      2867: begin
        W_PARAM = 16116;
      end
      2868: begin
        W_PARAM = 16019;
      end
      2869: begin
        W_PARAM = 16099;
      end
      2870: begin
        W_PARAM = 48778;
      end
      2871: begin
        W_PARAM = 48860;
      end
      2872: begin
        W_PARAM = 48553;
      end
      2873: begin
        W_PARAM = 15919;
      end
      2874: begin
        W_PARAM = 48725;
      end
      2875: begin
        W_PARAM = 16125;
      end
      2876: begin
        W_PARAM = 15648;
      end
      2877: begin
        W_PARAM = 15896;
      end
      2878: begin
        W_PARAM = 15948;
      end
      2879: begin
        W_PARAM = 48502;
      end
      2880: begin
        W_PARAM = 48743;
      end
      2881: begin
        W_PARAM = 15785;
      end
      2882: begin
        W_PARAM = 15435;
      end
      2883: begin
        W_PARAM = 48789;
      end
      2884: begin
        W_PARAM = 48762;
      end
      2885: begin
        W_PARAM = 16179;
      end
      2886: begin
        W_PARAM = 15893;
      end
      2887: begin
        W_PARAM = 48654;
      end
      2888: begin
        W_PARAM = 15492;
      end
      2889: begin
        W_PARAM = 48482;
      end
      2890: begin
        W_PARAM = 16049;
      end
      2891: begin
        W_PARAM = 48851;
      end
      2892: begin
        W_PARAM = 48892;
      end
      2893: begin
        W_PARAM = 48978;
      end
      2894: begin
        W_PARAM = 15997;
      end
      2895: begin
        W_PARAM = 16145;
      end
      2896: begin
        W_PARAM = 48847;
      end
      2897: begin
        W_PARAM = 16104;
      end
      2898: begin
        W_PARAM = 16009;
      end
      2899: begin
        W_PARAM = 15996;
      end
      2900: begin
        W_PARAM = 48793;
      end
      2901: begin
        W_PARAM = 48253;
      end
      2902: begin
        W_PARAM = 16005;
      end
      2903: begin
        W_PARAM = 48843;
      end
      2904: begin
        W_PARAM = 48696;
      end
      2905: begin
        W_PARAM = 16041;
      end
      2906: begin
        W_PARAM = 48676;
      end
      2907: begin
        W_PARAM = 48545;
      end
      2908: begin
        W_PARAM = 16064;
      end
      2909: begin
        W_PARAM = 15912;
      end
      2910: begin
        W_PARAM = 16106;
      end
      2911: begin
        W_PARAM = 16081;
      end
      2912: begin
        W_PARAM = 16015;
      end
      2913: begin
        W_PARAM = 48862;
      end
      2914: begin
        W_PARAM = 48719;
      end
      2915: begin
        W_PARAM = 15911;
      end
      2916: begin
        W_PARAM = 48790;
      end
      2917: begin
        W_PARAM = 48893;
      end
      2918: begin
        W_PARAM = 16046;
      end
      2919: begin
        W_PARAM = 48744;
      end
      2920: begin
        W_PARAM = 48822;
      end
      2921: begin
        W_PARAM = 48771;
      end
      2922: begin
        W_PARAM = 16014;
      end
      2923: begin
        W_PARAM = 48965;
      end
      2924: begin
        W_PARAM = 16120;
      end
      2925: begin
        W_PARAM = 16128;
      end
      2926: begin
        W_PARAM = 48819;
      end
      2927: begin
        W_PARAM = 48881;
      end
      2928: begin
        W_PARAM = 16174;
      end
      2929: begin
        W_PARAM = 16004;
      end
      2930: begin
        W_PARAM = 16033;
      end
      2931: begin
        W_PARAM = 16144;
      end
      2932: begin
        W_PARAM = 48513;
      end
      2933: begin
        W_PARAM = 15873;
      end
      2934: begin
        W_PARAM = 48895;
      end
      2935: begin
        W_PARAM = 48243;
      end
      2936: begin
        W_PARAM = 48653;
      end
      2937: begin
        W_PARAM = 16048;
      end
      2938: begin
        W_PARAM = 15552;
      end
      2939: begin
        W_PARAM = 48937;
      end
      2940: begin
        W_PARAM = 16117;
      end
      2941: begin
        W_PARAM = 16117;
      end
      2942: begin
        W_PARAM = 16002;
      end
      2943: begin
        W_PARAM = 15880;
      end
      2944: begin
        W_PARAM = 49038;
      end
      2945: begin
        W_PARAM = 15412;
      end
      2946: begin
        W_PARAM = 48909;
      end
      2947: begin
        W_PARAM = 16086;
      end
      2948: begin
        W_PARAM = 48542;
      end
      2949: begin
        W_PARAM = 48387;
      end
      2950: begin
        W_PARAM = 48771;
      end
      2951: begin
        W_PARAM = 16260;
      end
      2952: begin
        W_PARAM = 48804;
      end
      2953: begin
        W_PARAM = 15522;
      end
      2954: begin
        W_PARAM = 15564;
      end
      2955: begin
        W_PARAM = 48506;
      end
      2956: begin
        W_PARAM = 48910;
      end
      2957: begin
        W_PARAM = 16189;
      end
      2958: begin
        W_PARAM = 48902;
      end
      2959: begin
        W_PARAM = 48580;
      end
      2960: begin
        W_PARAM = 16109;
      end
      2961: begin
        W_PARAM = 15992;
      end
      2962: begin
        W_PARAM = 48595;
      end
      2963: begin
        W_PARAM = 16026;
      end
      2964: begin
        W_PARAM = 48955;
      end
      2965: begin
        W_PARAM = 48815;
      end
      2966: begin
        W_PARAM = 48933;
      end
      2967: begin
        W_PARAM = 16283;
      end
      2968: begin
        W_PARAM = 48877;
      end
      2969: begin
        W_PARAM = 15756;
      end
      2970: begin
        W_PARAM = 16164;
      end
      2971: begin
        W_PARAM = 16020;
      end
      2972: begin
        W_PARAM = 16157;
      end
      2973: begin
        W_PARAM = 16030;
      end
      2974: begin
        W_PARAM = 47917;
      end
      2975: begin
        W_PARAM = 48926;
      end
      2976: begin
        W_PARAM = 48867;
      end
      2977: begin
        W_PARAM = 15410;
      end
      2978: begin
        W_PARAM = 48877;
      end
      2979: begin
        W_PARAM = 48812;
      end
      2980: begin
        W_PARAM = 16143;
      end
      2981: begin
        W_PARAM = 48811;
      end
      2982: begin
        W_PARAM = 15878;
      end
      2983: begin
        W_PARAM = 15891;
      end
      2984: begin
        W_PARAM = 48689;
      end
      2985: begin
        W_PARAM = 48942;
      end
      2986: begin
        W_PARAM = 48907;
      end
      2987: begin
        W_PARAM = 16025;
      end
      2988: begin
        W_PARAM = 16134;
      end
      2989: begin
        W_PARAM = 15766;
      end
      2990: begin
        W_PARAM = 48798;
      end
      2991: begin
        W_PARAM = 48401;
      end
      2992: begin
        W_PARAM = 48768;
      end
      2993: begin
        W_PARAM = 15873;
      end
      2994: begin
        W_PARAM = 16071;
      end
      2995: begin
        W_PARAM = 48907;
      end
      2996: begin
        W_PARAM = 48974;
      end
      2997: begin
        W_PARAM = 16147;
      end
      2998: begin
        W_PARAM = 16182;
      end
      2999: begin
        W_PARAM = 15890;
      end
      3000: begin
        W_PARAM = 15990;
      end
      3001: begin
        W_PARAM = 48951;
      end
      3002: begin
        W_PARAM = 48612;
      end
      3003: begin
        W_PARAM = 16119;
      end
      3004: begin
        W_PARAM = 48726;
      end
      3005: begin
        W_PARAM = 48829;
      end
      3006: begin
        W_PARAM = 48706;
      end
      3007: begin
        W_PARAM = 16180;
      end
      3008: begin
        W_PARAM = 15896;
      end
      3009: begin
        W_PARAM = 15522;
      end
      3010: begin
        W_PARAM = 15952;
      end
      3011: begin
        W_PARAM = 48531;
      end
      3012: begin
        W_PARAM = 48674;
      end
      3013: begin
        W_PARAM = 48790;
      end
      3014: begin
        W_PARAM = 15546;
      end
      3015: begin
        W_PARAM = 48400;
      end
      3016: begin
        W_PARAM = 48780;
      end
      3017: begin
        W_PARAM = 16093;
      end
      3018: begin
        W_PARAM = 16032;
      end
      3019: begin
        W_PARAM = 48653;
      end
      3020: begin
        W_PARAM = 16129;
      end
      3021: begin
        W_PARAM = 48899;
      end
      3022: begin
        W_PARAM = 48824;
      end
      3023: begin
        W_PARAM = 16008;
      end
      3024: begin
        W_PARAM = 15915;
      end
      3025: begin
        W_PARAM = 48825;
      end
      3026: begin
        W_PARAM = 48939;
      end
      3027: begin
        W_PARAM = 16054;
      end
      3028: begin
        W_PARAM = 16133;
      end
      3029: begin
        W_PARAM = 15799;
      end
      3030: begin
        W_PARAM = 16161;
      end
      3031: begin
        W_PARAM = 48939;
      end
      3032: begin
        W_PARAM = 48767;
      end
      3033: begin
        W_PARAM = 15983;
      end
      3034: begin
        W_PARAM = 48974;
      end
      3035: begin
        W_PARAM = 16224;
      end
      3036: begin
        W_PARAM = 15931;
      end
      3037: begin
        W_PARAM = 48830;
      end
      3038: begin
        W_PARAM = 16064;
      end
      3039: begin
        W_PARAM = 48722;
      end
      3040: begin
        W_PARAM = 16215;
      end
      3041: begin
        W_PARAM = 48953;
      end
      3042: begin
        W_PARAM = 49042;
      end
      3043: begin
        W_PARAM = 48987;
      end
      3044: begin
        W_PARAM = 48810;
      end
      3045: begin
        W_PARAM = 16450;
      end
      3046: begin
        W_PARAM = 15545;
      end
      3047: begin
        W_PARAM = 48672;
      end
      3048: begin
        W_PARAM = 48650;
      end
      3049: begin
        W_PARAM = 48912;
      end
      3050: begin
        W_PARAM = 48925;
      end
      3051: begin
        W_PARAM = 48773;
      end
      3052: begin
        W_PARAM = 48622;
      end
      3053: begin
        W_PARAM = 15593;
      end
      3054: begin
        W_PARAM = 48801;
      end
      3055: begin
        W_PARAM = 16398;
      end
      3056: begin
        W_PARAM = 49019;
      end
      3057: begin
        W_PARAM = 15926;
      end
      3058: begin
        W_PARAM = 48755;
      end
      3059: begin
        W_PARAM = 15820;
      end
      3060: begin
        W_PARAM = 48848;
      end
      3061: begin
        W_PARAM = 48542;
      end
      3062: begin
        W_PARAM = 15922;
      end
      3063: begin
        W_PARAM = 48212;
      end
      3064: begin
        W_PARAM = 48803;
      end
      3065: begin
        W_PARAM = 16227;
      end
      3066: begin
        W_PARAM = 48847;
      end
      3067: begin
        W_PARAM = 15836;
      end
      3068: begin
        W_PARAM = 15925;
      end
      3069: begin
        W_PARAM = 48644;
      end
      3070: begin
        W_PARAM = 47609;
      end
      3071: begin
        W_PARAM = 15416;
      end
      3072: begin
        W_PARAM = 47831;
      end
      3073: begin
        W_PARAM = 47394;
      end
      3074: begin
        W_PARAM = 48030;
      end
      3075: begin
        W_PARAM = 47954;
      end
      3076: begin
        W_PARAM = 48446;
      end
      3077: begin
        W_PARAM = 15770;
      end
      3078: begin
        W_PARAM = 48203;
      end
      3079: begin
        W_PARAM = 48270;
      end
      3080: begin
        W_PARAM = 46475;
      end
      3081: begin
        W_PARAM = 46919;
      end
      3082: begin
        W_PARAM = 47167;
      end
      3083: begin
        W_PARAM = 47644;
      end
      3084: begin
        W_PARAM = 47360;
      end
      3085: begin
        W_PARAM = 47121;
      end
      3086: begin
        W_PARAM = 45980;
      end
      3087: begin
        W_PARAM = 15042;
      end
      3088: begin
        W_PARAM = 46740;
      end
      3089: begin
        W_PARAM = 47661;
      end
      3090: begin
        W_PARAM = 15678;
      end
      3091: begin
        W_PARAM = 14987;
      end
      3092: begin
        W_PARAM = 47794;
      end
      3093: begin
        W_PARAM = 48345;
      end
      3094: begin
        W_PARAM = 48538;
      end
      3095: begin
        W_PARAM = 48338;
      end
      3096: begin
        W_PARAM = 47447;
      end
      3097: begin
        W_PARAM = 16008;
      end
      3098: begin
        W_PARAM = 47988;
      end
      3099: begin
        W_PARAM = 48697;
      end
      3100: begin
        W_PARAM = 47755;
      end
      3101: begin
        W_PARAM = 47265;
      end
      3102: begin
        W_PARAM = 48457;
      end
      3103: begin
        W_PARAM = 48148;
      end
      3104: begin
        W_PARAM = 48802;
      end
      3105: begin
        W_PARAM = 48470;
      end
      3106: begin
        W_PARAM = 47872;
      end
      3107: begin
        W_PARAM = 16271;
      end
      3108: begin
        W_PARAM = 48411;
      end
      3109: begin
        W_PARAM = 48935;
      end
      3110: begin
        W_PARAM = 15856;
      end
      3111: begin
        W_PARAM = 48640;
      end
      3112: begin
        W_PARAM = 48429;
      end
      3113: begin
        W_PARAM = 16254;
      end
      3114: begin
        W_PARAM = 15869;
      end
      3115: begin
        W_PARAM = 48996;
      end
      3116: begin
        W_PARAM = 48710;
      end
      3117: begin
        W_PARAM = 16057;
      end
      3118: begin
        W_PARAM = 15573;
      end
      3119: begin
        W_PARAM = 48828;
      end
      3120: begin
        W_PARAM = 48901;
      end
      3121: begin
        W_PARAM = 48726;
      end
      3122: begin
        W_PARAM = 48810;
      end
      3123: begin
        W_PARAM = 16210;
      end
      3124: begin
        W_PARAM = 48845;
      end
      3125: begin
        W_PARAM = 48632;
      end
      3126: begin
        W_PARAM = 15894;
      end
      3127: begin
        W_PARAM = 16160;
      end
      3128: begin
        W_PARAM = 15881;
      end
      3129: begin
        W_PARAM = 48657;
      end
      3130: begin
        W_PARAM = 48808;
      end
      3131: begin
        W_PARAM = 48828;
      end
      3132: begin
        W_PARAM = 16017;
      end
      3133: begin
        W_PARAM = 48716;
      end
      3134: begin
        W_PARAM = 15726;
      end
      3135: begin
        W_PARAM = 48664;
      end
      3136: begin
        W_PARAM = 16006;
      end
      3137: begin
        W_PARAM = 15429;
      end
      3138: begin
        W_PARAM = 16077;
      end
      3139: begin
        W_PARAM = 15561;
      end
      3140: begin
        W_PARAM = 15937;
      end
      3141: begin
        W_PARAM = 49044;
      end
      3142: begin
        W_PARAM = 16088;
      end
      3143: begin
        W_PARAM = 48775;
      end
      3144: begin
        W_PARAM = 16084;
      end
      3145: begin
        W_PARAM = 16061;
      end
      3146: begin
        W_PARAM = 48772;
      end
      3147: begin
        W_PARAM = 15691;
      end
      3148: begin
        W_PARAM = 15887;
      end
      3149: begin
        W_PARAM = 15807;
      end
      3150: begin
        W_PARAM = 15931;
      end
      3151: begin
        W_PARAM = 48961;
      end
      3152: begin
        W_PARAM = 15605;
      end
      3153: begin
        W_PARAM = 49005;
      end
      3154: begin
        W_PARAM = 48598;
      end
      3155: begin
        W_PARAM = 15909;
      end
      3156: begin
        W_PARAM = 16043;
      end
      3157: begin
        W_PARAM = 15891;
      end
      3158: begin
        W_PARAM = 16182;
      end
      3159: begin
        W_PARAM = 15975;
      end
      3160: begin
        W_PARAM = 15937;
      end
      3161: begin
        W_PARAM = 48874;
      end
      3162: begin
        W_PARAM = 48950;
      end
      3163: begin
        W_PARAM = 48672;
      end
      3164: begin
        W_PARAM = 15866;
      end
      3165: begin
        W_PARAM = 15897;
      end
      3166: begin
        W_PARAM = 48660;
      end
      3167: begin
        W_PARAM = 48917;
      end
      3168: begin
        W_PARAM = 16140;
      end
      3169: begin
        W_PARAM = 16262;
      end
      3170: begin
        W_PARAM = 48919;
      end
      3171: begin
        W_PARAM = 48934;
      end
      3172: begin
        W_PARAM = 48835;
      end
      3173: begin
        W_PARAM = 48917;
      end
      3174: begin
        W_PARAM = 16172;
      end
      3175: begin
        W_PARAM = 15872;
      end
      3176: begin
        W_PARAM = 16084;
      end
      3177: begin
        W_PARAM = 16040;
      end
      3178: begin
        W_PARAM = 16149;
      end
      3179: begin
        W_PARAM = 15772;
      end
      3180: begin
        W_PARAM = 48655;
      end
      3181: begin
        W_PARAM = 48850;
      end
      3182: begin
        W_PARAM = 49051;
      end
      3183: begin
        W_PARAM = 48920;
      end
      3184: begin
        W_PARAM = 16234;
      end
      3185: begin
        W_PARAM = 48455;
      end
      3186: begin
        W_PARAM = 48684;
      end
      3187: begin
        W_PARAM = 16200;
      end
      3188: begin
        W_PARAM = 16009;
      end
      3189: begin
        W_PARAM = 16155;
      end
      3190: begin
        W_PARAM = 15673;
      end
      3191: begin
        W_PARAM = 48470;
      end
      3192: begin
        W_PARAM = 48973;
      end
      3193: begin
        W_PARAM = 48735;
      end
      3194: begin
        W_PARAM = 48708;
      end
      3195: begin
        W_PARAM = 15954;
      end
      3196: begin
        W_PARAM = 48783;
      end
      3197: begin
        W_PARAM = 16128;
      end
      3198: begin
        W_PARAM = 16050;
      end
      3199: begin
        W_PARAM = 16099;
      end
      3200: begin
        W_PARAM = 49021;
      end
      3201: begin
        W_PARAM = 48855;
      end
      3202: begin
        W_PARAM = 49025;
      end
      3203: begin
        W_PARAM = 15610;
      end
      3204: begin
        W_PARAM = 16282;
      end
      3205: begin
        W_PARAM = 15876;
      end
      3206: begin
        W_PARAM = 16081;
      end
      3207: begin
        W_PARAM = 48312;
      end
      3208: begin
        W_PARAM = 15886;
      end
      3209: begin
        W_PARAM = 16136;
      end
      3210: begin
        W_PARAM = 48476;
      end
      3211: begin
        W_PARAM = 16167;
      end
      3212: begin
        W_PARAM = 49079;
      end
      3213: begin
        W_PARAM = 16100;
      end
      3214: begin
        W_PARAM = 49103;
      end
      3215: begin
        W_PARAM = 16213;
      end
      3216: begin
        W_PARAM = 16066;
      end
      3217: begin
        W_PARAM = 16007;
      end
      3218: begin
        W_PARAM = 16061;
      end
      3219: begin
        W_PARAM = 15914;
      end
      3220: begin
        W_PARAM = 48923;
      end
      3221: begin
        W_PARAM = 16178;
      end
      3222: begin
        W_PARAM = 48948;
      end
      3223: begin
        W_PARAM = 15472;
      end
      3224: begin
        W_PARAM = 49040;
      end
      3225: begin
        W_PARAM = 15765;
      end
      3226: begin
        W_PARAM = 48816;
      end
      3227: begin
        W_PARAM = 16208;
      end
      3228: begin
        W_PARAM = 16266;
      end
      3229: begin
        W_PARAM = 15831;
      end
      3230: begin
        W_PARAM = 49012;
      end
      3231: begin
        W_PARAM = 16256;
      end
      3232: begin
        W_PARAM = 48929;
      end
      3233: begin
        W_PARAM = 16051;
      end
      3234: begin
        W_PARAM = 16208;
      end
      3235: begin
        W_PARAM = 48809;
      end
      3236: begin
        W_PARAM = 49004;
      end
      3237: begin
        W_PARAM = 16035;
      end
      3238: begin
        W_PARAM = 48590;
      end
      3239: begin
        W_PARAM = 16105;
      end
      3240: begin
        W_PARAM = 49042;
      end
      3241: begin
        W_PARAM = 16022;
      end
      3242: begin
        W_PARAM = 48751;
      end
      3243: begin
        W_PARAM = 48785;
      end
      3244: begin
        W_PARAM = 16192;
      end
      3245: begin
        W_PARAM = 48815;
      end
      3246: begin
        W_PARAM = 15757;
      end
      3247: begin
        W_PARAM = 16122;
      end
      3248: begin
        W_PARAM = 48532;
      end
      3249: begin
        W_PARAM = 16115;
      end
      3250: begin
        W_PARAM = 15820;
      end
      3251: begin
        W_PARAM = 48777;
      end
      3252: begin
        W_PARAM = 48936;
      end
      3253: begin
        W_PARAM = 16152;
      end
      3254: begin
        W_PARAM = 16019;
      end
      3255: begin
        W_PARAM = 48775;
      end
      3256: begin
        W_PARAM = 48955;
      end
      3257: begin
        W_PARAM = 16107;
      end
      3258: begin
        W_PARAM = 48781;
      end
      3259: begin
        W_PARAM = 16193;
      end
      3260: begin
        W_PARAM = 48942;
      end
      3261: begin
        W_PARAM = 48152;
      end
      3262: begin
        W_PARAM = 15706;
      end
      3263: begin
        W_PARAM = 15959;
      end
      3264: begin
        W_PARAM = 15962;
      end
      3265: begin
        W_PARAM = 48441;
      end
      3266: begin
        W_PARAM = 48890;
      end
      3267: begin
        W_PARAM = 16169;
      end
      3268: begin
        W_PARAM = 48848;
      end
      3269: begin
        W_PARAM = 16125;
      end
      3270: begin
        W_PARAM = 15874;
      end
      3271: begin
        W_PARAM = 48777;
      end
      3272: begin
        W_PARAM = 16154;
      end
      3273: begin
        W_PARAM = 48408;
      end
      3274: begin
        W_PARAM = 15618;
      end
      3275: begin
        W_PARAM = 48910;
      end
      3276: begin
        W_PARAM = 48504;
      end
      3277: begin
        W_PARAM = 15723;
      end
      3278: begin
        W_PARAM = 48516;
      end
      3279: begin
        W_PARAM = 15915;
      end
      3280: begin
        W_PARAM = 15824;
      end
      3281: begin
        W_PARAM = 48617;
      end
      3282: begin
        W_PARAM = 48824;
      end
      3283: begin
        W_PARAM = 16098;
      end
      3284: begin
        W_PARAM = 48758;
      end
      3285: begin
        W_PARAM = 49032;
      end
      3286: begin
        W_PARAM = 48659;
      end
      3287: begin
        W_PARAM = 16147;
      end
      3288: begin
        W_PARAM = 48334;
      end
      3289: begin
        W_PARAM = 16212;
      end
      3290: begin
        W_PARAM = 16235;
      end
      3291: begin
        W_PARAM = 48807;
      end
      3292: begin
        W_PARAM = 15974;
      end
      3293: begin
        W_PARAM = 48615;
      end
      3294: begin
        W_PARAM = 48931;
      end
      3295: begin
        W_PARAM = 48921;
      end
      3296: begin
        W_PARAM = 48091;
      end
      3297: begin
        W_PARAM = 15963;
      end
      3298: begin
        W_PARAM = 48489;
      end
      3299: begin
        W_PARAM = 16065;
      end
      3300: begin
        W_PARAM = 16075;
      end
      3301: begin
        W_PARAM = 48840;
      end
      3302: begin
        W_PARAM = 48472;
      end
      3303: begin
        W_PARAM = 16048;
      end
      3304: begin
        W_PARAM = 48885;
      end
      3305: begin
        W_PARAM = 49037;
      end
      3306: begin
        W_PARAM = 48841;
      end
      3307: begin
        W_PARAM = 16191;
      end
      3308: begin
        W_PARAM = 16065;
      end
      3309: begin
        W_PARAM = 16142;
      end
      3310: begin
        W_PARAM = 15899;
      end
      3311: begin
        W_PARAM = 48825;
      end
      3312: begin
        W_PARAM = 48562;
      end
      3313: begin
        W_PARAM = 48750;
      end
      3314: begin
        W_PARAM = 49000;
      end
      3315: begin
        W_PARAM = 16211;
      end
      3316: begin
        W_PARAM = 16185;
      end
      3317: begin
        W_PARAM = 48807;
      end
      3318: begin
        W_PARAM = 16142;
      end
      3319: begin
        W_PARAM = 48816;
      end
      3320: begin
        W_PARAM = 16132;
      end
      3321: begin
        W_PARAM = 48904;
      end
      3322: begin
        W_PARAM = 48785;
      end
      3323: begin
        W_PARAM = 48948;
      end
      3324: begin
        W_PARAM = 49028;
      end
      3325: begin
        W_PARAM = 16390;
      end
      3326: begin
        W_PARAM = 15909;
      end
      3327: begin
        W_PARAM = 48812;
      end
      3328: begin
        W_PARAM = 16162;
      end
      3329: begin
        W_PARAM = 48901;
      end
      3330: begin
        W_PARAM = 48872;
      end
      3331: begin
        W_PARAM = 48800;
      end
      3332: begin
        W_PARAM = 15923;
      end
      3333: begin
        W_PARAM = 15897;
      end
      3334: begin
        W_PARAM = 48893;
      end
      3335: begin
        W_PARAM = 16417;
      end
      3336: begin
        W_PARAM = 49035;
      end
      3337: begin
        W_PARAM = 48771;
      end
      3338: begin
        W_PARAM = 48300;
      end
      3339: begin
        W_PARAM = 48735;
      end
      3340: begin
        W_PARAM = 48821;
      end
      3341: begin
        W_PARAM = 48577;
      end
      3342: begin
        W_PARAM = 15875;
      end
      3343: begin
        W_PARAM = 48012;
      end
      3344: begin
        W_PARAM = 48686;
      end
      3345: begin
        W_PARAM = 16194;
      end
      3346: begin
        W_PARAM = 48972;
      end
      3347: begin
        W_PARAM = 48311;
      end
      3348: begin
        W_PARAM = 16160;
      end
      3349: begin
        W_PARAM = 48526;
      end
      3350: begin
        W_PARAM = 47763;
      end
      3351: begin
        W_PARAM = 15625;
      end
      3352: begin
        W_PARAM = 48540;
      end
      3353: begin
        W_PARAM = 47377;
      end
      3354: begin
        W_PARAM = 47932;
      end
      3355: begin
        W_PARAM = 15271;
      end
      3356: begin
        W_PARAM = 15664;
      end
      3357: begin
        W_PARAM = 15512;
      end
      3358: begin
        W_PARAM = 48259;
      end
      3359: begin
        W_PARAM = 47985;
      end
      3360: begin
        W_PARAM = 46110;
      end
      3361: begin
        W_PARAM = 45315;
      end
      3362: begin
        W_PARAM = 47154;
      end
      3363: begin
        W_PARAM = 47601;
      end
      3364: begin
        W_PARAM = 46120;
      end
      3365: begin
        W_PARAM = 46899;
      end
      3366: begin
        W_PARAM = 44626;
      end
      3367: begin
        W_PARAM = 15136;
      end
      3368: begin
        W_PARAM = 46717;
      end
      3369: begin
        W_PARAM = 47869;
      end
      3370: begin
        W_PARAM = 14741;
      end
      3371: begin
        W_PARAM = 47412;
      end
      3372: begin
        W_PARAM = 47374;
      end
      3373: begin
        W_PARAM = 48176;
      end
      3374: begin
        W_PARAM = 48552;
      end
      3375: begin
        W_PARAM = 48424;
      end
      3376: begin
        W_PARAM = 47558;
      end
      3377: begin
        W_PARAM = 15966;
      end
      3378: begin
        W_PARAM = 47887;
      end
      3379: begin
        W_PARAM = 48548;
      end
      3380: begin
        W_PARAM = 47886;
      end
      3381: begin
        W_PARAM = 48281;
      end
      3382: begin
        W_PARAM = 47906;
      end
      3383: begin
        W_PARAM = 48424;
      end
      3384: begin
        W_PARAM = 48837;
      end
      3385: begin
        W_PARAM = 48468;
      end
      3386: begin
        W_PARAM = 47868;
      end
      3387: begin
        W_PARAM = 16260;
      end
      3388: begin
        W_PARAM = 48378;
      end
      3389: begin
        W_PARAM = 48895;
      end
      3390: begin
        W_PARAM = 48143;
      end
      3391: begin
        W_PARAM = 48171;
      end
      3392: begin
        W_PARAM = 48868;
      end
      3393: begin
        W_PARAM = 15920;
      end
      3394: begin
        W_PARAM = 48746;
      end
      3395: begin
        W_PARAM = 48804;
      end
      3396: begin
        W_PARAM = 48676;
      end
      3397: begin
        W_PARAM = 16229;
      end
      3398: begin
        W_PARAM = 16114;
      end
      3399: begin
        W_PARAM = 48829;
      end
      3400: begin
        W_PARAM = 48708;
      end
      3401: begin
        W_PARAM = 15787;
      end
      3402: begin
        W_PARAM = 48793;
      end
      3403: begin
        W_PARAM = 15316;
      end
      3404: begin
        W_PARAM = 48960;
      end
      3405: begin
        W_PARAM = 15340;
      end
      3406: begin
        W_PARAM = 15757;
      end
      3407: begin
        W_PARAM = 16229;
      end
      3408: begin
        W_PARAM = 48712;
      end
      3409: begin
        W_PARAM = 16065;
      end
      3410: begin
        W_PARAM = 15417;
      end
      3411: begin
        W_PARAM = 48652;
      end
      3412: begin
        W_PARAM = 48920;
      end
      3413: begin
        W_PARAM = 48764;
      end
      3414: begin
        W_PARAM = 15592;
      end
      3415: begin
        W_PARAM = 48644;
      end
      3416: begin
        W_PARAM = 48708;
      end
      3417: begin
        W_PARAM = 16069;
      end
      3418: begin
        W_PARAM = 16129;
      end
      3419: begin
        W_PARAM = 16061;
      end
      3420: begin
        W_PARAM = 16169;
      end
      3421: begin
        W_PARAM = 48761;
      end
      3422: begin
        W_PARAM = 49064;
      end
      3423: begin
        W_PARAM = 48896;
      end
      3424: begin
        W_PARAM = 15896;
      end
      3425: begin
        W_PARAM = 16197;
      end
      3426: begin
        W_PARAM = 15652;
      end
      3427: begin
        W_PARAM = 48672;
      end
      3428: begin
        W_PARAM = 48675;
      end
      3429: begin
        W_PARAM = 16192;
      end
      3430: begin
        W_PARAM = 48646;
      end
      3431: begin
        W_PARAM = 48819;
      end
      3432: begin
        W_PARAM = 49130;
      end
      3433: begin
        W_PARAM = 48773;
      end
      3434: begin
        W_PARAM = 16143;
      end
      3435: begin
        W_PARAM = 15852;
      end
      3436: begin
        W_PARAM = 16106;
      end
      3437: begin
        W_PARAM = 16194;
      end
      3438: begin
        W_PARAM = 16075;
      end
      3439: begin
        W_PARAM = 16013;
      end
      3440: begin
        W_PARAM = 48708;
      end
      3441: begin
        W_PARAM = 48862;
      end
      3442: begin
        W_PARAM = 48926;
      end
      3443: begin
        W_PARAM = 48972;
      end
      3444: begin
        W_PARAM = 16168;
      end
      3445: begin
        W_PARAM = 15746;
      end
      3446: begin
        W_PARAM = 16115;
      end
      3447: begin
        W_PARAM = 16257;
      end
      3448: begin
        W_PARAM = 48757;
      end
      3449: begin
        W_PARAM = 15772;
      end
      3450: begin
        W_PARAM = 48174;
      end
      3451: begin
        W_PARAM = 48566;
      end
      3452: begin
        W_PARAM = 48902;
      end
      3453: begin
        W_PARAM = 48654;
      end
      3454: begin
        W_PARAM = 15359;
      end
      3455: begin
        W_PARAM = 48808;
      end
      3456: begin
        W_PARAM = 16099;
      end
      3457: begin
        W_PARAM = 48692;
      end
      3458: begin
        W_PARAM = 15936;
      end
      3459: begin
        W_PARAM = 16160;
      end
      3460: begin
        W_PARAM = 48496;
      end
      3461: begin
        W_PARAM = 48878;
      end
      3462: begin
        W_PARAM = 48896;
      end
      3463: begin
        W_PARAM = 16128;
      end
      3464: begin
        W_PARAM = 16161;
      end
      3465: begin
        W_PARAM = 16104;
      end
      3466: begin
        W_PARAM = 48526;
      end
      3467: begin
        W_PARAM = 48863;
      end
      3468: begin
        W_PARAM = 48748;
      end
      3469: begin
        W_PARAM = 15927;
      end
      3470: begin
        W_PARAM = 15920;
      end
      3471: begin
        W_PARAM = 48930;
      end
      3472: begin
        W_PARAM = 49007;
      end
      3473: begin
        W_PARAM = 48843;
      end
      3474: begin
        W_PARAM = 16145;
      end
      3475: begin
        W_PARAM = 48267;
      end
      3476: begin
        W_PARAM = 16192;
      end
      3477: begin
        W_PARAM = 16037;
      end
      3478: begin
        W_PARAM = 48732;
      end
      3479: begin
        W_PARAM = 16069;
      end
      3480: begin
        W_PARAM = 16068;
      end
      3481: begin
        W_PARAM = 15928;
      end
      3482: begin
        W_PARAM = 48926;
      end
      3483: begin
        W_PARAM = 15511;
      end
      3484: begin
        W_PARAM = 16307;
      end
      3485: begin
        W_PARAM = 15759;
      end
      3486: begin
        W_PARAM = 48222;
      end
      3487: begin
        W_PARAM = 49021;
      end
      3488: begin
        W_PARAM = 15934;
      end
      3489: begin
        W_PARAM = 48924;
      end
      3490: begin
        W_PARAM = 16009;
      end
      3491: begin
        W_PARAM = 15814;
      end
      3492: begin
        W_PARAM = 48759;
      end
      3493: begin
        W_PARAM = 48779;
      end
      3494: begin
        W_PARAM = 16072;
      end
      3495: begin
        W_PARAM = 16083;
      end
      3496: begin
        W_PARAM = 16018;
      end
      3497: begin
        W_PARAM = 49117;
      end
      3498: begin
        W_PARAM = 16164;
      end
      3499: begin
        W_PARAM = 15898;
      end
      3500: begin
        W_PARAM = 48934;
      end
      3501: begin
        W_PARAM = 16292;
      end
      3502: begin
        W_PARAM = 48955;
      end
      3503: begin
        W_PARAM = 16200;
      end
      3504: begin
        W_PARAM = 49004;
      end
      3505: begin
        W_PARAM = 48739;
      end
      3506: begin
        W_PARAM = 48775;
      end
      3507: begin
        W_PARAM = 15884;
      end
      3508: begin
        W_PARAM = 15971;
      end
      3509: begin
        W_PARAM = 16060;
      end
      3510: begin
        W_PARAM = 49041;
      end
      3511: begin
        W_PARAM = 16083;
      end
      3512: begin
        W_PARAM = 48934;
      end
      3513: begin
        W_PARAM = 15931;
      end
      3514: begin
        W_PARAM = 48518;
      end
      3515: begin
        W_PARAM = 16016;
      end
      3516: begin
        W_PARAM = 48849;
      end
      3517: begin
        W_PARAM = 16193;
      end
      3518: begin
        W_PARAM = 15736;
      end
      3519: begin
        W_PARAM = 16143;
      end
      3520: begin
        W_PARAM = 48946;
      end
      3521: begin
        W_PARAM = 16088;
      end
      3522: begin
        W_PARAM = 48734;
      end
      3523: begin
        W_PARAM = 16001;
      end
      3524: begin
        W_PARAM = 16066;
      end
      3525: begin
        W_PARAM = 48884;
      end
      3526: begin
        W_PARAM = 48787;
      end
      3527: begin
        W_PARAM = 16115;
      end
      3528: begin
        W_PARAM = 48576;
      end
      3529: begin
        W_PARAM = 15994;
      end
      3530: begin
        W_PARAM = 15841;
      end
      3531: begin
        W_PARAM = 15812;
      end
      3532: begin
        W_PARAM = 48821;
      end
      3533: begin
        W_PARAM = 48789;
      end
      3534: begin
        W_PARAM = 48465;
      end
      3535: begin
        W_PARAM = 48948;
      end
      3536: begin
        W_PARAM = 48408;
      end
      3537: begin
        W_PARAM = 16161;
      end
      3538: begin
        W_PARAM = 16035;
      end
      3539: begin
        W_PARAM = 16016;
      end
      3540: begin
        W_PARAM = 48700;
      end
      3541: begin
        W_PARAM = 48726;
      end
      3542: begin
        W_PARAM = 48893;
      end
      3543: begin
        W_PARAM = 15904;
      end
      3544: begin
        W_PARAM = 48382;
      end
      3545: begin
        W_PARAM = 48832;
      end
      3546: begin
        W_PARAM = 48713;
      end
      3547: begin
        W_PARAM = 16171;
      end
      3548: begin
        W_PARAM = 48431;
      end
      3549: begin
        W_PARAM = 16181;
      end
      3550: begin
        W_PARAM = 16039;
      end
      3551: begin
        W_PARAM = 48838;
      end
      3552: begin
        W_PARAM = 16072;
      end
      3553: begin
        W_PARAM = 48787;
      end
      3554: begin
        W_PARAM = 16000;
      end
      3555: begin
        W_PARAM = 48920;
      end
      3556: begin
        W_PARAM = 48953;
      end
      3557: begin
        W_PARAM = 48598;
      end
      3558: begin
        W_PARAM = 16162;
      end
      3559: begin
        W_PARAM = 16123;
      end
      3560: begin
        W_PARAM = 15944;
      end
      3561: begin
        W_PARAM = 48678;
      end
      3562: begin
        W_PARAM = 15758;
      end
      3563: begin
        W_PARAM = 16012;
      end
      3564: begin
        W_PARAM = 15891;
      end
      3565: begin
        W_PARAM = 48792;
      end
      3566: begin
        W_PARAM = 48806;
      end
      3567: begin
        W_PARAM = 48780;
      end
      3568: begin
        W_PARAM = 15945;
      end
      3569: begin
        W_PARAM = 15927;
      end
      3570: begin
        W_PARAM = 15743;
      end
      3571: begin
        W_PARAM = 48309;
      end
      3572: begin
        W_PARAM = 48514;
      end
      3573: begin
        W_PARAM = 49025;
      end
      3574: begin
        W_PARAM = 16192;
      end
      3575: begin
        W_PARAM = 49066;
      end
      3576: begin
        W_PARAM = 15737;
      end
      3577: begin
        W_PARAM = 15828;
      end
      3578: begin
        W_PARAM = 16199;
      end
      3579: begin
        W_PARAM = 16170;
      end
      3580: begin
        W_PARAM = 16011;
      end
      3581: begin
        W_PARAM = 48487;
      end
      3582: begin
        W_PARAM = 15660;
      end
      3583: begin
        W_PARAM = 48970;
      end
      3584: begin
        W_PARAM = 15970;
      end
      3585: begin
        W_PARAM = 49155;
      end
      3586: begin
        W_PARAM = 16191;
      end
      3587: begin
        W_PARAM = 16126;
      end
      3588: begin
        W_PARAM = 16064;
      end
      3589: begin
        W_PARAM = 16188;
      end
      3590: begin
        W_PARAM = 16100;
      end
      3591: begin
        W_PARAM = 48371;
      end
      3592: begin
        W_PARAM = 48983;
      end
      3593: begin
        W_PARAM = 48919;
      end
      3594: begin
        W_PARAM = 48441;
      end
      3595: begin
        W_PARAM = 49171;
      end
      3596: begin
        W_PARAM = 16301;
      end
      3597: begin
        W_PARAM = 48889;
      end
      3598: begin
        W_PARAM = 16297;
      end
      3599: begin
        W_PARAM = 16277;
      end
      3600: begin
        W_PARAM = 16305;
      end
      3601: begin
        W_PARAM = 48669;
      end
      3602: begin
        W_PARAM = 16150;
      end
      3603: begin
        W_PARAM = 48807;
      end
      3604: begin
        W_PARAM = 15809;
      end
      3605: begin
        W_PARAM = 49211;
      end
      3606: begin
        W_PARAM = 16183;
      end
      3607: begin
        W_PARAM = 48896;
      end
      3608: begin
        W_PARAM = 16376;
      end
      3609: begin
        W_PARAM = 48979;
      end
      3610: begin
        W_PARAM = 48476;
      end
      3611: begin
        W_PARAM = 48608;
      end
      3612: begin
        W_PARAM = 16184;
      end
      3613: begin
        W_PARAM = 15886;
      end
      3614: begin
        W_PARAM = 48680;
      end
      3615: begin
        W_PARAM = 15875;
      end
      3616: begin
        W_PARAM = 48819;
      end
      3617: begin
        W_PARAM = 15761;
      end
      3618: begin
        W_PARAM = 15604;
      end
      3619: begin
        W_PARAM = 48849;
      end
      3620: begin
        W_PARAM = 48807;
      end
      3621: begin
        W_PARAM = 48642;
      end
      3622: begin
        W_PARAM = 16171;
      end
      3623: begin
        W_PARAM = 47705;
      end
      3624: begin
        W_PARAM = 48663;
      end
      3625: begin
        W_PARAM = 16216;
      end
      3626: begin
        W_PARAM = 48998;
      end
      3627: begin
        W_PARAM = 15941;
      end
      3628: begin
        W_PARAM = 48522;
      end
      3629: begin
        W_PARAM = 48650;
      end
      3630: begin
        W_PARAM = 47873;
      end
      3631: begin
        W_PARAM = 15591;
      end
      3632: begin
        W_PARAM = 15524;
      end
      3633: begin
        W_PARAM = 47492;
      end
      3634: begin
        W_PARAM = 48443;
      end
      3635: begin
        W_PARAM = 48286;
      end
      3636: begin
        W_PARAM = 15513;
      end
      3637: begin
        W_PARAM = 15788;
      end
      3638: begin
        W_PARAM = 48545;
      end
      3639: begin
        W_PARAM = 48038;
      end
      3640: begin
        W_PARAM = 45039;
      end
      3641: begin
        W_PARAM = 14532;
      end
      3642: begin
        W_PARAM = 46899;
      end
      3643: begin
        W_PARAM = 47122;
      end
      3644: begin
        W_PARAM = 45981;
      end
      3645: begin
        W_PARAM = 46475;
      end
      3646: begin
        W_PARAM = 46346;
      end
      3647: begin
        W_PARAM = 47036;
      end
      3648: begin
        W_PARAM = 46746;
      end
      3649: begin
        W_PARAM = 47009;
      end
      3650: begin
        W_PARAM = 15000;
      end
      3651: begin
        W_PARAM = 47086;
      end
      3652: begin
        W_PARAM = 47204;
      end
      3653: begin
        W_PARAM = 47862;
      end
      3654: begin
        W_PARAM = 48519;
      end
      3655: begin
        W_PARAM = 48076;
      end
      3656: begin
        W_PARAM = 47606;
      end
      3657: begin
        W_PARAM = 15859;
      end
      3658: begin
        W_PARAM = 47476;
      end
      3659: begin
        W_PARAM = 48441;
      end
      3660: begin
        W_PARAM = 48046;
      end
      3661: begin
        W_PARAM = 48061;
      end
      3662: begin
        W_PARAM = 47682;
      end
      3663: begin
        W_PARAM = 48211;
      end
      3664: begin
        W_PARAM = 48783;
      end
      3665: begin
        W_PARAM = 48249;
      end
      3666: begin
        W_PARAM = 47407;
      end
      3667: begin
        W_PARAM = 16169;
      end
      3668: begin
        W_PARAM = 48095;
      end
      3669: begin
        W_PARAM = 48811;
      end
      3670: begin
        W_PARAM = 48278;
      end
      3671: begin
        W_PARAM = 15752;
      end
      3672: begin
        W_PARAM = 48918;
      end
      3673: begin
        W_PARAM = 15910;
      end
      3674: begin
        W_PARAM = 48788;
      end
      3675: begin
        W_PARAM = 15648;
      end
      3676: begin
        W_PARAM = 48656;
      end
      3677: begin
        W_PARAM = 16220;
      end
      3678: begin
        W_PARAM = 16034;
      end
      3679: begin
        W_PARAM = 48849;
      end
      3680: begin
        W_PARAM = 16072;
      end
      3681: begin
        W_PARAM = 15989;
      end
      3682: begin
        W_PARAM = 49109;
      end
      3683: begin
        W_PARAM = 48938;
      end
      3684: begin
        W_PARAM = 48757;
      end
      3685: begin
        W_PARAM = 16012;
      end
      3686: begin
        W_PARAM = 15646;
      end
      3687: begin
        W_PARAM = 16103;
      end
      3688: begin
        W_PARAM = 48815;
      end
      3689: begin
        W_PARAM = 16322;
      end
      3690: begin
        W_PARAM = 48776;
      end
      3691: begin
        W_PARAM = 48595;
      end
      3692: begin
        W_PARAM = 49071;
      end
      3693: begin
        W_PARAM = 48716;
      end
      3694: begin
        W_PARAM = 16005;
      end
      3695: begin
        W_PARAM = 16147;
      end
      3696: begin
        W_PARAM = 15986;
      end
      3697: begin
        W_PARAM = 15724;
      end
      3698: begin
        W_PARAM = 15967;
      end
      3699: begin
        W_PARAM = 16152;
      end
      3700: begin
        W_PARAM = 16152;
      end
      3701: begin
        W_PARAM = 48681;
      end
      3702: begin
        W_PARAM = 49112;
      end
      3703: begin
        W_PARAM = 48792;
      end
      3704: begin
        W_PARAM = 16169;
      end
      3705: begin
        W_PARAM = 48913;
      end
      3706: begin
        W_PARAM = 16232;
      end
      3707: begin
        W_PARAM = 16157;
      end
      3708: begin
        W_PARAM = 48437;
      end
      3709: begin
        W_PARAM = 48302;
      end
      3710: begin
        W_PARAM = 16075;
      end
      3711: begin
        W_PARAM = 48822;
      end
      3712: begin
        W_PARAM = 49047;
      end
      3713: begin
        W_PARAM = 48849;
      end
      3714: begin
        W_PARAM = 16056;
      end
      3715: begin
        W_PARAM = 16057;
      end
      3716: begin
        W_PARAM = 15626;
      end
      3717: begin
        W_PARAM = 15780;
      end
      3718: begin
        W_PARAM = 15893;
      end
      3719: begin
        W_PARAM = 16146;
      end
      3720: begin
        W_PARAM = 15705;
      end
      3721: begin
        W_PARAM = 15932;
      end
      3722: begin
        W_PARAM = 48819;
      end
      3723: begin
        W_PARAM = 48676;
      end
      3724: begin
        W_PARAM = 16100;
      end
      3725: begin
        W_PARAM = 48640;
      end
      3726: begin
        W_PARAM = 48658;
      end
      3727: begin
        W_PARAM = 48775;
      end
      3728: begin
        W_PARAM = 48309;
      end
      3729: begin
        W_PARAM = 16067;
      end
      3730: begin
        W_PARAM = 15746;
      end
      3731: begin
        W_PARAM = 16009;
      end
      3732: begin
        W_PARAM = 48882;
      end
      3733: begin
        W_PARAM = 48676;
      end
      3734: begin
        W_PARAM = 16152;
      end
      3735: begin
        W_PARAM = 15793;
      end
      3736: begin
        W_PARAM = 48636;
      end
      3737: begin
        W_PARAM = 48778;
      end
      3738: begin
        W_PARAM = 15992;
      end
      3739: begin
        W_PARAM = 48746;
      end
      3740: begin
        W_PARAM = 16132;
      end
      3741: begin
        W_PARAM = 49017;
      end
      3742: begin
        W_PARAM = 48893;
      end
      3743: begin
        W_PARAM = 48811;
      end
      3744: begin
        W_PARAM = 16200;
      end
      3745: begin
        W_PARAM = 15946;
      end
      3746: begin
        W_PARAM = 16091;
      end
      3747: begin
        W_PARAM = 15737;
      end
      3748: begin
        W_PARAM = 48806;
      end
      3749: begin
        W_PARAM = 15890;
      end
      3750: begin
        W_PARAM = 48283;
      end
      3751: begin
        W_PARAM = 49009;
      end
      3752: begin
        W_PARAM = 16014;
      end
      3753: begin
        W_PARAM = 48694;
      end
      3754: begin
        W_PARAM = 16212;
      end
      3755: begin
        W_PARAM = 16003;
      end
      3756: begin
        W_PARAM = 48908;
      end
      3757: begin
        W_PARAM = 15806;
      end
      3758: begin
        W_PARAM = 15939;
      end
      3759: begin
        W_PARAM = 15645;
      end
      3760: begin
        W_PARAM = 15631;
      end
      3761: begin
        W_PARAM = 16081;
      end
      3762: begin
        W_PARAM = 48770;
      end
      3763: begin
        W_PARAM = 15905;
      end
      3764: begin
        W_PARAM = 16130;
      end
      3765: begin
        W_PARAM = 16198;
      end
      3766: begin
        W_PARAM = 15929;
      end
      3767: begin
        W_PARAM = 49105;
      end
      3768: begin
        W_PARAM = 15993;
      end
      3769: begin
        W_PARAM = 48854;
      end
      3770: begin
        W_PARAM = 49036;
      end
      3771: begin
        W_PARAM = 16096;
      end
      3772: begin
        W_PARAM = 16045;
      end
      3773: begin
        W_PARAM = 16117;
      end
      3774: begin
        W_PARAM = 48905;
      end
      3775: begin
        W_PARAM = 16065;
      end
      3776: begin
        W_PARAM = 16106;
      end
      3777: begin
        W_PARAM = 49086;
      end
      3778: begin
        W_PARAM = 16222;
      end
      3779: begin
        W_PARAM = 15908;
      end
      3780: begin
        W_PARAM = 48983;
      end
      3781: begin
        W_PARAM = 16105;
      end
      3782: begin
        W_PARAM = 15773;
      end
      3783: begin
        W_PARAM = 16038;
      end
      3784: begin
        W_PARAM = 16010;
      end
      3785: begin
        W_PARAM = 48783;
      end
      3786: begin
        W_PARAM = 48806;
      end
      3787: begin
        W_PARAM = 15954;
      end
      3788: begin
        W_PARAM = 48803;
      end
      3789: begin
        W_PARAM = 16093;
      end
      3790: begin
        W_PARAM = 49049;
      end
      3791: begin
        W_PARAM = 16089;
      end
      3792: begin
        W_PARAM = 48835;
      end
      3793: begin
        W_PARAM = 48856;
      end
      3794: begin
        W_PARAM = 16191;
      end
      3795: begin
        W_PARAM = 48833;
      end
      3796: begin
        W_PARAM = 15645;
      end
      3797: begin
        W_PARAM = 15512;
      end
      3798: begin
        W_PARAM = 16185;
      end
      3799: begin
        W_PARAM = 16092;
      end
      3800: begin
        W_PARAM = 48942;
      end
      3801: begin
        W_PARAM = 15531;
      end
      3802: begin
        W_PARAM = 48891;
      end
      3803: begin
        W_PARAM = 15904;
      end
      3804: begin
        W_PARAM = 16022;
      end
      3805: begin
        W_PARAM = 48914;
      end
      3806: begin
        W_PARAM = 15593;
      end
      3807: begin
        W_PARAM = 16074;
      end
      3808: begin
        W_PARAM = 15795;
      end
      3809: begin
        W_PARAM = 16195;
      end
      3810: begin
        W_PARAM = 48833;
      end
      3811: begin
        W_PARAM = 16231;
      end
      3812: begin
        W_PARAM = 48501;
      end
      3813: begin
        W_PARAM = 15766;
      end
      3814: begin
        W_PARAM = 15798;
      end
      3815: begin
        W_PARAM = 48669;
      end
      3816: begin
        W_PARAM = 48880;
      end
      3817: begin
        W_PARAM = 48603;
      end
      3818: begin
        W_PARAM = 48672;
      end
      3819: begin
        W_PARAM = 16002;
      end
      3820: begin
        W_PARAM = 15730;
      end
      3821: begin
        W_PARAM = 48823;
      end
      3822: begin
        W_PARAM = 48824;
      end
      3823: begin
        W_PARAM = 16022;
      end
      3824: begin
        W_PARAM = 16059;
      end
      3825: begin
        W_PARAM = 48560;
      end
      3826: begin
        W_PARAM = 48755;
      end
      3827: begin
        W_PARAM = 48466;
      end
      3828: begin
        W_PARAM = 15771;
      end
      3829: begin
        W_PARAM = 16024;
      end
      3830: begin
        W_PARAM = 15766;
      end
      3831: begin
        W_PARAM = 48906;
      end
      3832: begin
        W_PARAM = 48840;
      end
      3833: begin
        W_PARAM = 16029;
      end
      3834: begin
        W_PARAM = 48404;
      end
      3835: begin
        W_PARAM = 16022;
      end
      3836: begin
        W_PARAM = 16025;
      end
      3837: begin
        W_PARAM = 48932;
      end
      3838: begin
        W_PARAM = 48535;
      end
      3839: begin
        W_PARAM = 16181;
      end
      3840: begin
        W_PARAM = 48949;
      end
      3841: begin
        W_PARAM = 48675;
      end
      3842: begin
        W_PARAM = 48886;
      end
      3843: begin
        W_PARAM = 48957;
      end
      3844: begin
        W_PARAM = 16125;
      end
      3845: begin
        W_PARAM = 48405;
      end
      3846: begin
        W_PARAM = 48772;
      end
      3847: begin
        W_PARAM = 16140;
      end
      3848: begin
        W_PARAM = 16176;
      end
      3849: begin
        W_PARAM = 16167;
      end
      3850: begin
        W_PARAM = 48836;
      end
      3851: begin
        W_PARAM = 48702;
      end
      3852: begin
        W_PARAM = 15684;
      end
      3853: begin
        W_PARAM = 48938;
      end
      3854: begin
        W_PARAM = 16143;
      end
      3855: begin
        W_PARAM = 48794;
      end
      3856: begin
        W_PARAM = 16183;
      end
      3857: begin
        W_PARAM = 16132;
      end
      3858: begin
        W_PARAM = 48916;
      end
      3859: begin
        W_PARAM = 16011;
      end
      3860: begin
        W_PARAM = 16051;
      end
      3861: begin
        W_PARAM = 48787;
      end
      3862: begin
        W_PARAM = 15821;
      end
      3863: begin
        W_PARAM = 49085;
      end
      3864: begin
        W_PARAM = 16140;
      end
      3865: begin
        W_PARAM = 15379;
      end
      3866: begin
        W_PARAM = 16011;
      end
      3867: begin
        W_PARAM = 48731;
      end
      3868: begin
        W_PARAM = 15982;
      end
      3869: begin
        W_PARAM = 16115;
      end
      3870: begin
        W_PARAM = 16143;
      end
      3871: begin
        W_PARAM = 48776;
      end
      3872: begin
        W_PARAM = 48737;
      end
      3873: begin
        W_PARAM = 48890;
      end
      3874: begin
        W_PARAM = 48568;
      end
      3875: begin
        W_PARAM = 49019;
      end
      3876: begin
        W_PARAM = 16297;
      end
      3877: begin
        W_PARAM = 48815;
      end
      3878: begin
        W_PARAM = 16232;
      end
      3879: begin
        W_PARAM = 48841;
      end
      3880: begin
        W_PARAM = 16190;
      end
      3881: begin
        W_PARAM = 48801;
      end
      3882: begin
        W_PARAM = 16335;
      end
      3883: begin
        W_PARAM = 48653;
      end
      3884: begin
        W_PARAM = 48930;
      end
      3885: begin
        W_PARAM = 49155;
      end
      3886: begin
        W_PARAM = 16224;
      end
      3887: begin
        W_PARAM = 15963;
      end
      3888: begin
        W_PARAM = 16212;
      end
      3889: begin
        W_PARAM = 49043;
      end
      3890: begin
        W_PARAM = 16136;
      end
      3891: begin
        W_PARAM = 48744;
      end
      3892: begin
        W_PARAM = 16315;
      end
      3893: begin
        W_PARAM = 15758;
      end
      3894: begin
        W_PARAM = 15954;
      end
      3895: begin
        W_PARAM = 49000;
      end
      3896: begin
        W_PARAM = 48939;
      end
      3897: begin
        W_PARAM = 15943;
      end
      3898: begin
        W_PARAM = 48079;
      end
      3899: begin
        W_PARAM = 48935;
      end
      3900: begin
        W_PARAM = 48560;
      end
      3901: begin
        W_PARAM = 48647;
      end
      3902: begin
        W_PARAM = 16331;
      end
      3903: begin
        W_PARAM = 47943;
      end
      3904: begin
        W_PARAM = 48541;
      end
      3905: begin
        W_PARAM = 48479;
      end
      3906: begin
        W_PARAM = 48979;
      end
      3907: begin
        W_PARAM = 15539;
      end
      3908: begin
        W_PARAM = 48731;
      end
      3909: begin
        W_PARAM = 48734;
      end
      3910: begin
        W_PARAM = 48180;
      end
      3911: begin
        W_PARAM = 47757;
      end
      3912: begin
        W_PARAM = 16155;
      end
      3913: begin
        W_PARAM = 48235;
      end
      3914: begin
        W_PARAM = 48688;
      end
      3915: begin
        W_PARAM = 48694;
      end
      3916: begin
        W_PARAM = 48672;
      end
      3917: begin
        W_PARAM = 48492;
      end
      3918: begin
        W_PARAM = 48239;
      end
      3919: begin
        W_PARAM = 47947;
      end
      3920: begin
        W_PARAM = 46979;
      end
      3921: begin
        W_PARAM = 46440;
      end
      3922: begin
        W_PARAM = 47172;
      end
      3923: begin
        W_PARAM = 48075;
      end
      3924: begin
        W_PARAM = 47496;
      end
      3925: begin
        W_PARAM = 15618;
      end
      3926: begin
        W_PARAM = 47549;
      end
      3927: begin
        W_PARAM = 47327;
      end
      3928: begin
        W_PARAM = 47578;
      end
      3929: begin
        W_PARAM = 48326;
      end
      3930: begin
        W_PARAM = 46992;
      end
      3931: begin
        W_PARAM = 46826;
      end
      3932: begin
        W_PARAM = 48511;
      end
      3933: begin
        W_PARAM = 15747;
      end
      3934: begin
        W_PARAM = 48425;
      end
      3935: begin
        W_PARAM = 47923;
      end
      3936: begin
        W_PARAM = 46854;
      end
      3937: begin
        W_PARAM = 15759;
      end
      3938: begin
        W_PARAM = 47655;
      end
      3939: begin
        W_PARAM = 48346;
      end
      3940: begin
        W_PARAM = 48070;
      end
      3941: begin
        W_PARAM = 15368;
      end
      3942: begin
        W_PARAM = 48421;
      end
      3943: begin
        W_PARAM = 15641;
      end
      3944: begin
        W_PARAM = 48630;
      end
      3945: begin
        W_PARAM = 48112;
      end
      3946: begin
        W_PARAM = 46954;
      end
      3947: begin
        W_PARAM = 16066;
      end
      3948: begin
        W_PARAM = 47886;
      end
      3949: begin
        W_PARAM = 48766;
      end
      3950: begin
        W_PARAM = 48843;
      end
      3951: begin
        W_PARAM = 15875;
      end
      3952: begin
        W_PARAM = 48895;
      end
      3953: begin
        W_PARAM = 15948;
      end
      3954: begin
        W_PARAM = 48404;
      end
      3955: begin
        W_PARAM = 15929;
      end
      3956: begin
        W_PARAM = 48527;
      end
      3957: begin
        W_PARAM = 16099;
      end
      3958: begin
        W_PARAM = 15601;
      end
      3959: begin
        W_PARAM = 15527;
      end
      3960: begin
        W_PARAM = 48739;
      end
      3961: begin
        W_PARAM = 15951;
      end
      3962: begin
        W_PARAM = 49007;
      end
      3963: begin
        W_PARAM = 48825;
      end
      3964: begin
        W_PARAM = 16274;
      end
      3965: begin
        W_PARAM = 16008;
      end
      3966: begin
        W_PARAM = 48927;
      end
      3967: begin
        W_PARAM = 16091;
      end
      3968: begin
        W_PARAM = 48913;
      end
      3969: begin
        W_PARAM = 16171;
      end
      3970: begin
        W_PARAM = 16056;
      end
      3971: begin
        W_PARAM = 48660;
      end
      3972: begin
        W_PARAM = 49056;
      end
      3973: begin
        W_PARAM = 48981;
      end
      3974: begin
        W_PARAM = 16223;
      end
      3975: begin
        W_PARAM = 48424;
      end
      3976: begin
        W_PARAM = 15969;
      end
      3977: begin
        W_PARAM = 16065;
      end
      3978: begin
        W_PARAM = 16107;
      end
      3979: begin
        W_PARAM = 48298;
      end
      3980: begin
        W_PARAM = 15367;
      end
      3981: begin
        W_PARAM = 48772;
      end
      3982: begin
        W_PARAM = 48577;
      end
      3983: begin
        W_PARAM = 48970;
      end
      3984: begin
        W_PARAM = 16032;
      end
      3985: begin
        W_PARAM = 48604;
      end
      3986: begin
        W_PARAM = 16059;
      end
      3987: begin
        W_PARAM = 48784;
      end
      3988: begin
        W_PARAM = 15907;
      end
      3989: begin
        W_PARAM = 16174;
      end
      3990: begin
        W_PARAM = 16243;
      end
      3991: begin
        W_PARAM = 48872;
      end
      3992: begin
        W_PARAM = 16165;
      end
      3993: begin
        W_PARAM = 48894;
      end
      3994: begin
        W_PARAM = 16168;
      end
      3995: begin
        W_PARAM = 48460;
      end
      3996: begin
        W_PARAM = 48713;
      end
      3997: begin
        W_PARAM = 48250;
      end
      3998: begin
        W_PARAM = 49041;
      end
      3999: begin
        W_PARAM = 15804;
      end
      4000: begin
        W_PARAM = 15873;
      end
      4001: begin
        W_PARAM = 15984;
      end
      4002: begin
        W_PARAM = 48702;
      end
      4003: begin
        W_PARAM = 48620;
      end
      4004: begin
        W_PARAM = 16059;
      end
      4005: begin
        W_PARAM = 15837;
      end
      4006: begin
        W_PARAM = 15904;
      end
      4007: begin
        W_PARAM = 48455;
      end
      4008: begin
        W_PARAM = 48902;
      end
      4009: begin
        W_PARAM = 48619;
      end
      4010: begin
        W_PARAM = 16141;
      end
      4011: begin
        W_PARAM = 48773;
      end
      4012: begin
        W_PARAM = 48768;
      end
      4013: begin
        W_PARAM = 48644;
      end
      4014: begin
        W_PARAM = 15958;
      end
      4015: begin
        W_PARAM = 15957;
      end
      4016: begin
        W_PARAM = 16168;
      end
      4017: begin
        W_PARAM = 48860;
      end
      4018: begin
        W_PARAM = 48921;
      end
      4019: begin
        W_PARAM = 15669;
      end
      4020: begin
        W_PARAM = 48920;
      end
      4021: begin
        W_PARAM = 48984;
      end
      4022: begin
        W_PARAM = 16006;
      end
      4023: begin
        W_PARAM = 48583;
      end
      4024: begin
        W_PARAM = 15986;
      end
      4025: begin
        W_PARAM = 16104;
      end
      4026: begin
        W_PARAM = 16142;
      end
      4027: begin
        W_PARAM = 48676;
      end
      4028: begin
        W_PARAM = 15855;
      end
      4029: begin
        W_PARAM = 15772;
      end
      4030: begin
        W_PARAM = 15941;
      end
      4031: begin
        W_PARAM = 48987;
      end
      4032: begin
        W_PARAM = 15942;
      end
      4033: begin
        W_PARAM = 48861;
      end
      4034: begin
        W_PARAM = 16069;
      end
      4035: begin
        W_PARAM = 48358;
      end
      4036: begin
        W_PARAM = 16209;
      end
      4037: begin
        W_PARAM = 48956;
      end
      4038: begin
        W_PARAM = 16093;
      end
      4039: begin
        W_PARAM = 15625;
      end
      4040: begin
        W_PARAM = 16187;
      end
      4041: begin
        W_PARAM = 15788;
      end
      4042: begin
        W_PARAM = 48702;
      end
      4043: begin
        W_PARAM = 16027;
      end
      4044: begin
        W_PARAM = 16154;
      end
      4045: begin
        W_PARAM = 15755;
      end
      4046: begin
        W_PARAM = 15688;
      end
      4047: begin
        W_PARAM = 49109;
      end
      4048: begin
        W_PARAM = 16008;
      end
      4049: begin
        W_PARAM = 48767;
      end
      4050: begin
        W_PARAM = 48625;
      end
      4051: begin
        W_PARAM = 15866;
      end
      4052: begin
        W_PARAM = 15953;
      end
      4053: begin
        W_PARAM = 48688;
      end
      4054: begin
        W_PARAM = 48840;
      end
      4055: begin
        W_PARAM = 48568;
      end
      4056: begin
        W_PARAM = 48471;
      end
      4057: begin
        W_PARAM = 48852;
      end
      4058: begin
        W_PARAM = 16162;
      end
      4059: begin
        W_PARAM = 16014;
      end
      4060: begin
        W_PARAM = 49059;
      end
      4061: begin
        W_PARAM = 16194;
      end
      4062: begin
        W_PARAM = 15858;
      end
      4063: begin
        W_PARAM = 15997;
      end
      4064: begin
        W_PARAM = 16010;
      end
      4065: begin
        W_PARAM = 15547;
      end
      4066: begin
        W_PARAM = 48860;
      end
      4067: begin
        W_PARAM = 48736;
      end
      4068: begin
        W_PARAM = 16014;
      end
      4069: begin
        W_PARAM = 15977;
      end
      4070: begin
        W_PARAM = 48928;
      end
      4071: begin
        W_PARAM = 16180;
      end
      4072: begin
        W_PARAM = 48841;
      end
      4073: begin
        W_PARAM = 15783;
      end
      4074: begin
        W_PARAM = 15827;
      end
      4075: begin
        W_PARAM = 48689;
      end
      4076: begin
        W_PARAM = 15607;
      end
      4077: begin
        W_PARAM = 48703;
      end
      4078: begin
        W_PARAM = 15942;
      end
      4079: begin
        W_PARAM = 16009;
      end
      4080: begin
        W_PARAM = 49073;
      end
      4081: begin
        W_PARAM = 16013;
      end
      4082: begin
        W_PARAM = 15499;
      end
      4083: begin
        W_PARAM = 48597;
      end
      4084: begin
        W_PARAM = 16136;
      end
      4085: begin
        W_PARAM = 48860;
      end
      4086: begin
        W_PARAM = 16144;
      end
      4087: begin
        W_PARAM = 15950;
      end
      4088: begin
        W_PARAM = 48608;
      end
      4089: begin
        W_PARAM = 16094;
      end
      4090: begin
        W_PARAM = 15788;
      end
      4091: begin
        W_PARAM = 48311;
      end
      4092: begin
        W_PARAM = 48914;
      end
      4093: begin
        W_PARAM = 15820;
      end
      4094: begin
        W_PARAM = 16167;
      end
      4095: begin
        W_PARAM = 48905;
      end
      4096: begin
        W_PARAM = 48983;
      end
      4097: begin
        W_PARAM = 16132;
      end
      4098: begin
        W_PARAM = 15915;
      end
      4099: begin
        W_PARAM = 16104;
      end
      4100: begin
        W_PARAM = 48494;
      end
      4101: begin
        W_PARAM = 49027;
      end
      4102: begin
        W_PARAM = 16129;
      end
      4103: begin
        W_PARAM = 15637;
      end
      4104: begin
        W_PARAM = 15920;
      end
      4105: begin
        W_PARAM = 48811;
      end
      4106: begin
        W_PARAM = 15537;
      end
      4107: begin
        W_PARAM = 16166;
      end
      4108: begin
        W_PARAM = 48786;
      end
      4109: begin
        W_PARAM = 16035;
      end
      4110: begin
        W_PARAM = 48784;
      end
      4111: begin
        W_PARAM = 48935;
      end
      4112: begin
        W_PARAM = 48746;
      end
      4113: begin
        W_PARAM = 48876;
      end
      4114: begin
        W_PARAM = 16187;
      end
      4115: begin
        W_PARAM = 48925;
      end
      4116: begin
        W_PARAM = 15793;
      end
      4117: begin
        W_PARAM = 16305;
      end
      4118: begin
        W_PARAM = 15751;
      end
      4119: begin
        W_PARAM = 48380;
      end
      4120: begin
        W_PARAM = 16025;
      end
      4121: begin
        W_PARAM = 48783;
      end
      4122: begin
        W_PARAM = 16067;
      end
      4123: begin
        W_PARAM = 48933;
      end
      4124: begin
        W_PARAM = 16047;
      end
      4125: begin
        W_PARAM = 15905;
      end
      4126: begin
        W_PARAM = 48862;
      end
      4127: begin
        W_PARAM = 16089;
      end
      4128: begin
        W_PARAM = 48878;
      end
      4129: begin
        W_PARAM = 15970;
      end
      4130: begin
        W_PARAM = 16157;
      end
      4131: begin
        W_PARAM = 48808;
      end
      4132: begin
        W_PARAM = 48797;
      end
      4133: begin
        W_PARAM = 16008;
      end
      4134: begin
        W_PARAM = 48538;
      end
      4135: begin
        W_PARAM = 48691;
      end
      4136: begin
        W_PARAM = 16005;
      end
      4137: begin
        W_PARAM = 48831;
      end
      4138: begin
        W_PARAM = 15756;
      end
      4139: begin
        W_PARAM = 15700;
      end
      4140: begin
        W_PARAM = 15912;
      end
      4141: begin
        W_PARAM = 48706;
      end
      4142: begin
        W_PARAM = 48447;
      end
      4143: begin
        W_PARAM = 48822;
      end
      4144: begin
        W_PARAM = 15972;
      end
      4145: begin
        W_PARAM = 16082;
      end
      4146: begin
        W_PARAM = 16049;
      end
      4147: begin
        W_PARAM = 16044;
      end
      4148: begin
        W_PARAM = 49003;
      end
      4149: begin
        W_PARAM = 15606;
      end
      4150: begin
        W_PARAM = 16133;
      end
      4151: begin
        W_PARAM = 48630;
      end
      4152: begin
        W_PARAM = 16133;
      end
      4153: begin
        W_PARAM = 48717;
      end
      4154: begin
        W_PARAM = 48744;
      end
      4155: begin
        W_PARAM = 16138;
      end
      4156: begin
        W_PARAM = 16053;
      end
      4157: begin
        W_PARAM = 16172;
      end
      4158: begin
        W_PARAM = 49027;
      end
      4159: begin
        W_PARAM = 49028;
      end
      4160: begin
        W_PARAM = 16244;
      end
      4161: begin
        W_PARAM = 48480;
      end
      4162: begin
        W_PARAM = 16060;
      end
      4163: begin
        W_PARAM = 15918;
      end
      4164: begin
        W_PARAM = 48904;
      end
      4165: begin
        W_PARAM = 16049;
      end
      4166: begin
        W_PARAM = 16184;
      end
      4167: begin
        W_PARAM = 48703;
      end
      4168: begin
        W_PARAM = 48908;
      end
      4169: begin
        W_PARAM = 49054;
      end
      4170: begin
        W_PARAM = 16099;
      end
      4171: begin
        W_PARAM = 48567;
      end
      4172: begin
        W_PARAM = 16250;
      end
      4173: begin
        W_PARAM = 48499;
      end
      4174: begin
        W_PARAM = 48505;
      end
      4175: begin
        W_PARAM = 49038;
      end
      4176: begin
        W_PARAM = 15892;
      end
      4177: begin
        W_PARAM = 48867;
      end
      4178: begin
        W_PARAM = 16135;
      end
      4179: begin
        W_PARAM = 48810;
      end
      4180: begin
        W_PARAM = 48392;
      end
      4181: begin
        W_PARAM = 48227;
      end
      4182: begin
        W_PARAM = 16274;
      end
      4183: begin
        W_PARAM = 48437;
      end
      4184: begin
        W_PARAM = 48831;
      end
      4185: begin
        W_PARAM = 48634;
      end
      4186: begin
        W_PARAM = 48893;
      end
      4187: begin
        W_PARAM = 48386;
      end
      4188: begin
        W_PARAM = 15368;
      end
      4189: begin
        W_PARAM = 48402;
      end
      4190: begin
        W_PARAM = 47609;
      end
      4191: begin
        W_PARAM = 47195;
      end
      4192: begin
        W_PARAM = 15718;
      end
      4193: begin
        W_PARAM = 48165;
      end
      4194: begin
        W_PARAM = 48282;
      end
      4195: begin
        W_PARAM = 48051;
      end
      4196: begin
        W_PARAM = 48281;
      end
      4197: begin
        W_PARAM = 47668;
      end
      4198: begin
        W_PARAM = 47858;
      end
      4199: begin
        W_PARAM = 47162;
      end
      4200: begin
        W_PARAM = 46775;
      end
      4201: begin
        W_PARAM = 46235;
      end
      4202: begin
        W_PARAM = 46977;
      end
      4203: begin
        W_PARAM = 47877;
      end
      4204: begin
        W_PARAM = 47291;
      end
      4205: begin
        W_PARAM = 15398;
      end
      4206: begin
        W_PARAM = 47351;
      end
      4207: begin
        W_PARAM = 14754;
      end
      4208: begin
        W_PARAM = 47377;
      end
      4209: begin
        W_PARAM = 48132;
      end
      4210: begin
        W_PARAM = 46850;
      end
      4211: begin
        W_PARAM = 46276;
      end
      4212: begin
        W_PARAM = 48646;
      end
      4213: begin
        W_PARAM = 15882;
      end
      4214: begin
        W_PARAM = 46477;
      end
      4215: begin
        W_PARAM = 47927;
      end
      4216: begin
        W_PARAM = 46087;
      end
      4217: begin
        W_PARAM = 46436;
      end
      4218: begin
        W_PARAM = 47779;
      end
      4219: begin
        W_PARAM = 46647;
      end
      4220: begin
        W_PARAM = 48044;
      end
      4221: begin
        W_PARAM = 15693;
      end
      4222: begin
        W_PARAM = 48543;
      end
      4223: begin
        W_PARAM = 15886;
      end
      4224: begin
        W_PARAM = 15830;
      end
      4225: begin
        W_PARAM = 48301;
      end
      4226: begin
        W_PARAM = 47535;
      end
      4227: begin
        W_PARAM = 15708;
      end
      4228: begin
        W_PARAM = 47906;
      end
      4229: begin
        W_PARAM = 48757;
      end
      4230: begin
        W_PARAM = 48867;
      end
      4231: begin
        W_PARAM = 15470;
      end
      4232: begin
        W_PARAM = 15691;
      end
      4233: begin
        W_PARAM = 15595;
      end
      4234: begin
        W_PARAM = 15986;
      end
      4235: begin
        W_PARAM = 48579;
      end
      4236: begin
        W_PARAM = 48700;
      end
      4237: begin
        W_PARAM = 16029;
      end
      4238: begin
        W_PARAM = 15318;
      end
      4239: begin
        W_PARAM = 15778;
      end
      4240: begin
        W_PARAM = 16085;
      end
      4241: begin
        W_PARAM = 15374;
      end
      4242: begin
        W_PARAM = 16053;
      end
      4243: begin
        W_PARAM = 15811;
      end
      4244: begin
        W_PARAM = 16134;
      end
      4245: begin
        W_PARAM = 47631;
      end
      4246: begin
        W_PARAM = 49033;
      end
      4247: begin
        W_PARAM = 48360;
      end
      4248: begin
        W_PARAM = 48870;
      end
      4249: begin
        W_PARAM = 15899;
      end
      4250: begin
        W_PARAM = 16153;
      end
      4251: begin
        W_PARAM = 48797;
      end
      4252: begin
        W_PARAM = 16268;
      end
      4253: begin
        W_PARAM = 48437;
      end
      4254: begin
        W_PARAM = 16022;
      end
      4255: begin
        W_PARAM = 48896;
      end
      4256: begin
        W_PARAM = 48851;
      end
      4257: begin
        W_PARAM = 48582;
      end
      4258: begin
        W_PARAM = 48951;
      end
      4259: begin
        W_PARAM = 15798;
      end
      4260: begin
        W_PARAM = 48945;
      end
      4261: begin
        W_PARAM = 48865;
      end
      4262: begin
        W_PARAM = 16144;
      end
      4263: begin
        W_PARAM = 16071;
      end
      4264: begin
        W_PARAM = 16129;
      end
      4265: begin
        W_PARAM = 15616;
      end
      4266: begin
        W_PARAM = 15927;
      end
      4267: begin
        W_PARAM = 48689;
      end
      4268: begin
        W_PARAM = 48898;
      end
      4269: begin
        W_PARAM = 15898;
      end
      4270: begin
        W_PARAM = 16168;
      end
      4271: begin
        W_PARAM = 48640;
      end
      4272: begin
        W_PARAM = 48912;
      end
      4273: begin
        W_PARAM = 48878;
      end
      4274: begin
        W_PARAM = 16146;
      end
      4275: begin
        W_PARAM = 48772;
      end
      4276: begin
        W_PARAM = 16111;
      end
      4277: begin
        W_PARAM = 48766;
      end
      4278: begin
        W_PARAM = 48701;
      end
      4279: begin
        W_PARAM = 15897;
      end
      4280: begin
        W_PARAM = 16042;
      end
      4281: begin
        W_PARAM = 15917;
      end
      4282: begin
        W_PARAM = 48662;
      end
      4283: begin
        W_PARAM = 48863;
      end
      4284: begin
        W_PARAM = 16023;
      end
      4285: begin
        W_PARAM = 15699;
      end
      4286: begin
        W_PARAM = 16029;
      end
      4287: begin
        W_PARAM = 48905;
      end
      4288: begin
        W_PARAM = 48752;
      end
      4289: begin
        W_PARAM = 15943;
      end
      4290: begin
        W_PARAM = 16085;
      end
      4291: begin
        W_PARAM = 48905;
      end
      4292: begin
        W_PARAM = 15965;
      end
      4293: begin
        W_PARAM = 48921;
      end
      4294: begin
        W_PARAM = 16128;
      end
      4295: begin
        W_PARAM = 16094;
      end
      4296: begin
        W_PARAM = 15266;
      end
      4297: begin
        W_PARAM = 48918;
      end
      4298: begin
        W_PARAM = 15913;
      end
      4299: begin
        W_PARAM = 48232;
      end
      4300: begin
        W_PARAM = 16194;
      end
      4301: begin
        W_PARAM = 48960;
      end
      4302: begin
        W_PARAM = 15426;
      end
      4303: begin
        W_PARAM = 48848;
      end
      4304: begin
        W_PARAM = 16139;
      end
      4305: begin
        W_PARAM = 48569;
      end
      4306: begin
        W_PARAM = 15889;
      end
      4307: begin
        W_PARAM = 47777;
      end
      4308: begin
        W_PARAM = 48814;
      end
      4309: begin
        W_PARAM = 15884;
      end
      4310: begin
        W_PARAM = 48648;
      end
      4311: begin
        W_PARAM = 15676;
      end
      4312: begin
        W_PARAM = 48424;
      end
      4313: begin
        W_PARAM = 48586;
      end
      4314: begin
        W_PARAM = 16136;
      end
      4315: begin
        W_PARAM = 15786;
      end
      4316: begin
        W_PARAM = 15973;
      end
      4317: begin
        W_PARAM = 48928;
      end
      4318: begin
        W_PARAM = 48631;
      end
      4319: begin
        W_PARAM = 15880;
      end
      4320: begin
        W_PARAM = 48639;
      end
      4321: begin
        W_PARAM = 16173;
      end
      4322: begin
        W_PARAM = 48582;
      end
      4323: begin
        W_PARAM = 15946;
      end
      4324: begin
        W_PARAM = 15830;
      end
      4325: begin
        W_PARAM = 15952;
      end
      4326: begin
        W_PARAM = 16114;
      end
      4327: begin
        W_PARAM = 49049;
      end
      4328: begin
        W_PARAM = 15833;
      end
      4329: begin
        W_PARAM = 48814;
      end
      4330: begin
        W_PARAM = 48964;
      end
      4331: begin
        W_PARAM = 16137;
      end
      4332: begin
        W_PARAM = 15986;
      end
      4333: begin
        W_PARAM = 48703;
      end
      4334: begin
        W_PARAM = 48860;
      end
      4335: begin
        W_PARAM = 47942;
      end
      4336: begin
        W_PARAM = 16054;
      end
      4337: begin
        W_PARAM = 48666;
      end
      4338: begin
        W_PARAM = 16079;
      end
      4339: begin
        W_PARAM = 15281;
      end
      4340: begin
        W_PARAM = 49074;
      end
      4341: begin
        W_PARAM = 16248;
      end
      4342: begin
        W_PARAM = 15908;
      end
      4343: begin
        W_PARAM = 16044;
      end
      4344: begin
        W_PARAM = 15899;
      end
      4345: begin
        W_PARAM = 48841;
      end
      4346: begin
        W_PARAM = 16123;
      end
      4347: begin
        W_PARAM = 48924;
      end
      4348: begin
        W_PARAM = 16177;
      end
      4349: begin
        W_PARAM = 48847;
      end
      4350: begin
        W_PARAM = 48939;
      end
      4351: begin
        W_PARAM = 48700;
      end
      4352: begin
        W_PARAM = 15852;
      end
      4353: begin
        W_PARAM = 15894;
      end
      4354: begin
        W_PARAM = 15934;
      end
      4355: begin
        W_PARAM = 48836;
      end
      4356: begin
        W_PARAM = 48711;
      end
      4357: begin
        W_PARAM = 16143;
      end
      4358: begin
        W_PARAM = 48530;
      end
      4359: begin
        W_PARAM = 16125;
      end
      4360: begin
        W_PARAM = 48925;
      end
      4361: begin
        W_PARAM = 16203;
      end
      4362: begin
        W_PARAM = 15593;
      end
      4363: begin
        W_PARAM = 15752;
      end
      4364: begin
        W_PARAM = 16171;
      end
      4365: begin
        W_PARAM = 48454;
      end
      4366: begin
        W_PARAM = 48707;
      end
      4367: begin
        W_PARAM = 48964;
      end
      4368: begin
        W_PARAM = 48604;
      end
      4369: begin
        W_PARAM = 15916;
      end
      4370: begin
        W_PARAM = 48892;
      end
      4371: begin
        W_PARAM = 48968;
      end
      4372: begin
        W_PARAM = 48858;
      end
      4373: begin
        W_PARAM = 48218;
      end
      4374: begin
        W_PARAM = 16182;
      end
      4375: begin
        W_PARAM = 48850;
      end
      4376: begin
        W_PARAM = 15861;
      end
      4377: begin
        W_PARAM = 16265;
      end
      4378: begin
        W_PARAM = 48847;
      end
      4379: begin
        W_PARAM = 16160;
      end
      4380: begin
        W_PARAM = 15795;
      end
      4381: begin
        W_PARAM = 48991;
      end
      4382: begin
        W_PARAM = 48797;
      end
      4383: begin
        W_PARAM = 48781;
      end
      4384: begin
        W_PARAM = 15768;
      end
      4385: begin
        W_PARAM = 16207;
      end
      4386: begin
        W_PARAM = 48594;
      end
      4387: begin
        W_PARAM = 16158;
      end
      4388: begin
        W_PARAM = 48310;
      end
      4389: begin
        W_PARAM = 48150;
      end
      4390: begin
        W_PARAM = 48050;
      end
      4391: begin
        W_PARAM = 49026;
      end
      4392: begin
        W_PARAM = 15935;
      end
      4393: begin
        W_PARAM = 15796;
      end
      4394: begin
        W_PARAM = 16109;
      end
      4395: begin
        W_PARAM = 15889;
      end
      4396: begin
        W_PARAM = 48533;
      end
      4397: begin
        W_PARAM = 48350;
      end
      4398: begin
        W_PARAM = 15304;
      end
      4399: begin
        W_PARAM = 15983;
      end
      4400: begin
        W_PARAM = 16076;
      end
      4401: begin
        W_PARAM = 48954;
      end
      4402: begin
        W_PARAM = 48929;
      end
      4403: begin
        W_PARAM = 16225;
      end
      4404: begin
        W_PARAM = 48836;
      end
      4405: begin
        W_PARAM = 48696;
      end
      4406: begin
        W_PARAM = 15856;
      end
      4407: begin
        W_PARAM = 16160;
      end
      4408: begin
        W_PARAM = 48666;
      end
      4409: begin
        W_PARAM = 15693;
      end
      4410: begin
        W_PARAM = 48456;
      end
      4411: begin
        W_PARAM = 48805;
      end
      4412: begin
        W_PARAM = 48531;
      end
      4413: begin
        W_PARAM = 16081;
      end
      4414: begin
        W_PARAM = 48841;
      end
      4415: begin
        W_PARAM = 15784;
      end
      4416: begin
        W_PARAM = 16052;
      end
      4417: begin
        W_PARAM = 16037;
      end
      4418: begin
        W_PARAM = 48609;
      end
      4419: begin
        W_PARAM = 48735;
      end
      4420: begin
        W_PARAM = 47676;
      end
      4421: begin
        W_PARAM = 48790;
      end
      4422: begin
        W_PARAM = 48983;
      end
      4423: begin
        W_PARAM = 16009;
      end
      4424: begin
        W_PARAM = 16219;
      end
      4425: begin
        W_PARAM = 48931;
      end
      4426: begin
        W_PARAM = 48791;
      end
      4427: begin
        W_PARAM = 16237;
      end
      4428: begin
        W_PARAM = 15883;
      end
      4429: begin
        W_PARAM = 48638;
      end
      4430: begin
        W_PARAM = 16094;
      end
      4431: begin
        W_PARAM = 48695;
      end
      4432: begin
        W_PARAM = 48876;
      end
      4433: begin
        W_PARAM = 16210;
      end
      4434: begin
        W_PARAM = 48555;
      end
      4435: begin
        W_PARAM = 15879;
      end
      4436: begin
        W_PARAM = 15621;
      end
      4437: begin
        W_PARAM = 16103;
      end
      4438: begin
        W_PARAM = 48921;
      end
      4439: begin
        W_PARAM = 48909;
      end
      4440: begin
        W_PARAM = 16253;
      end
      4441: begin
        W_PARAM = 48550;
      end
      4442: begin
        W_PARAM = 16269;
      end
      4443: begin
        W_PARAM = 16142;
      end
      4444: begin
        W_PARAM = 49078;
      end
      4445: begin
        W_PARAM = 16271;
      end
      4446: begin
        W_PARAM = 16043;
      end
      4447: begin
        W_PARAM = 48851;
      end
      4448: begin
        W_PARAM = 49026;
      end
      4449: begin
        W_PARAM = 49045;
      end
      4450: begin
        W_PARAM = 15891;
      end
      4451: begin
        W_PARAM = 48523;
      end
      4452: begin
        W_PARAM = 16244;
      end
      4453: begin
        W_PARAM = 48784;
      end
      4454: begin
        W_PARAM = 48777;
      end
      4455: begin
        W_PARAM = 48858;
      end
      4456: begin
        W_PARAM = 16213;
      end
      4457: begin
        W_PARAM = 48994;
      end
      4458: begin
        W_PARAM = 16077;
      end
      4459: begin
        W_PARAM = 48848;
      end
      4460: begin
        W_PARAM = 48474;
      end
      4461: begin
        W_PARAM = 48345;
      end
      4462: begin
        W_PARAM = 16257;
      end
      4463: begin
        W_PARAM = 48413;
      end
      4464: begin
        W_PARAM = 16003;
      end
      4465: begin
        W_PARAM = 48699;
      end
      4466: begin
        W_PARAM = 48907;
      end
      4467: begin
        W_PARAM = 48739;
      end
      4468: begin
        W_PARAM = 48434;
      end
      4469: begin
        W_PARAM = 48673;
      end
      4470: begin
        W_PARAM = 48044;
      end
      4471: begin
        W_PARAM = 47952;
      end
      4472: begin
        W_PARAM = 15970;
      end
      4473: begin
        W_PARAM = 47720;
      end
      4474: begin
        W_PARAM = 48420;
      end
      4475: begin
        W_PARAM = 48580;
      end
      4476: begin
        W_PARAM = 48494;
      end
      4477: begin
        W_PARAM = 47755;
      end
      4478: begin
        W_PARAM = 48002;
      end
      4479: begin
        W_PARAM = 48198;
      end
      4480: begin
        W_PARAM = 46596;
      end
      4481: begin
        W_PARAM = 45852;
      end
      4482: begin
        W_PARAM = 45711;
      end
      4483: begin
        W_PARAM = 46697;
      end
      4484: begin
        W_PARAM = 47054;
      end
      4485: begin
        W_PARAM = 47792;
      end
      4486: begin
        W_PARAM = 45561;
      end
      4487: begin
        W_PARAM = 15105;
      end
      4488: begin
        W_PARAM = 46880;
      end
      4489: begin
        W_PARAM = 47642;
      end
      4490: begin
        W_PARAM = 47272;
      end
      4491: begin
        W_PARAM = 14602;
      end
      4492: begin
        W_PARAM = 48513;
      end
      4493: begin
        W_PARAM = 15759;
      end
      4494: begin
        W_PARAM = 46446;
      end
      4495: begin
        W_PARAM = 47813;
      end
      4496: begin
        W_PARAM = 46604;
      end
      4497: begin
        W_PARAM = 47876;
      end
      4498: begin
        W_PARAM = 47921;
      end
      4499: begin
        W_PARAM = 47665;
      end
      4500: begin
        W_PARAM = 48263;
      end
      4501: begin
        W_PARAM = 15642;
      end
      4502: begin
        W_PARAM = 48351;
      end
      4503: begin
        W_PARAM = 16022;
      end
      4504: begin
        W_PARAM = 48212;
      end
      4505: begin
        W_PARAM = 48612;
      end
      4506: begin
        W_PARAM = 47871;
      end
      4507: begin
        W_PARAM = 48426;
      end
      4508: begin
        W_PARAM = 48146;
      end
      4509: begin
        W_PARAM = 48608;
      end
      4510: begin
        W_PARAM = 48771;
      end
      4511: begin
        W_PARAM = 47787;
      end
      4512: begin
        W_PARAM = 16262;
      end
      4513: begin
        W_PARAM = 15907;
      end
      4514: begin
        W_PARAM = 48727;
      end
      4515: begin
        W_PARAM = 48332;
      end
      4516: begin
        W_PARAM = 48777;
      end
      4517: begin
        W_PARAM = 48819;
      end
      4518: begin
        W_PARAM = 15687;
      end
      4519: begin
        W_PARAM = 48661;
      end
      4520: begin
        W_PARAM = 16150;
      end
      4521: begin
        W_PARAM = 48239;
      end
      4522: begin
        W_PARAM = 16197;
      end
      4523: begin
        W_PARAM = 16247;
      end
      4524: begin
        W_PARAM = 48988;
      end
      4525: begin
        W_PARAM = 48158;
      end
      4526: begin
        W_PARAM = 48998;
      end
      4527: begin
        W_PARAM = 48786;
      end
      4528: begin
        W_PARAM = 48882;
      end
      4529: begin
        W_PARAM = 15970;
      end
      4530: begin
        W_PARAM = 16179;
      end
      4531: begin
        W_PARAM = 48785;
      end
      4532: begin
        W_PARAM = 48456;
      end
      4533: begin
        W_PARAM = 16143;
      end
      4534: begin
        W_PARAM = 48820;
      end
      4535: begin
        W_PARAM = 15528;
      end
      4536: begin
        W_PARAM = 16060;
      end
      4537: begin
        W_PARAM = 48839;
      end
      4538: begin
        W_PARAM = 48954;
      end
      4539: begin
        W_PARAM = 15900;
      end
      4540: begin
        W_PARAM = 16102;
      end
      4541: begin
        W_PARAM = 48911;
      end
      4542: begin
        W_PARAM = 16157;
      end
      4543: begin
        W_PARAM = 48798;
      end
      4544: begin
        W_PARAM = 47753;
      end
      4545: begin
        W_PARAM = 48606;
      end
      4546: begin
        W_PARAM = 16142;
      end
      4547: begin
        W_PARAM = 48664;
      end
      4548: begin
        W_PARAM = 48633;
      end
      4549: begin
        W_PARAM = 48829;
      end
      4550: begin
        W_PARAM = 48362;
      end
      4551: begin
        W_PARAM = 48756;
      end
      4552: begin
        W_PARAM = 16023;
      end
      4553: begin
        W_PARAM = 48873;
      end
      4554: begin
        W_PARAM = 16122;
      end
      4555: begin
        W_PARAM = 49009;
      end
      4556: begin
        W_PARAM = 16148;
      end
      4557: begin
        W_PARAM = 16135;
      end
      4558: begin
        W_PARAM = 15755;
      end
      4559: begin
        W_PARAM = 48788;
      end
      4560: begin
        W_PARAM = 16147;
      end
      4561: begin
        W_PARAM = 48588;
      end
      4562: begin
        W_PARAM = 48846;
      end
      4563: begin
        W_PARAM = 48988;
      end
      4564: begin
        W_PARAM = 16134;
      end
      4565: begin
        W_PARAM = 48789;
      end
      4566: begin
        W_PARAM = 16044;
      end
      4567: begin
        W_PARAM = 48639;
      end
      4568: begin
        W_PARAM = 48404;
      end
      4569: begin
        W_PARAM = 16066;
      end
      4570: begin
        W_PARAM = 16086;
      end
      4571: begin
        W_PARAM = 16024;
      end
      4572: begin
        W_PARAM = 16030;
      end
      4573: begin
        W_PARAM = 15919;
      end
      4574: begin
        W_PARAM = 15845;
      end
      4575: begin
        W_PARAM = 48986;
      end
      4576: begin
        W_PARAM = 16115;
      end
      4577: begin
        W_PARAM = 48754;
      end
      4578: begin
        W_PARAM = 48534;
      end
      4579: begin
        W_PARAM = 48927;
      end
      4580: begin
        W_PARAM = 15886;
      end
      4581: begin
        W_PARAM = 48779;
      end
      4582: begin
        W_PARAM = 15932;
      end
      4583: begin
        W_PARAM = 48593;
      end
      4584: begin
        W_PARAM = 48774;
      end
      4585: begin
        W_PARAM = 15777;
      end
      4586: begin
        W_PARAM = 15988;
      end
      4587: begin
        W_PARAM = 48923;
      end
      4588: begin
        W_PARAM = 16114;
      end
      4589: begin
        W_PARAM = 15874;
      end
      4590: begin
        W_PARAM = 15950;
      end
      4591: begin
        W_PARAM = 48634;
      end
      4592: begin
        W_PARAM = 16033;
      end
      4593: begin
        W_PARAM = 48258;
      end
      4594: begin
        W_PARAM = 48663;
      end
      4595: begin
        W_PARAM = 48696;
      end
      4596: begin
        W_PARAM = 16293;
      end
      4597: begin
        W_PARAM = 49084;
      end
      4598: begin
        W_PARAM = 48030;
      end
      4599: begin
        W_PARAM = 15884;
      end
      4600: begin
        W_PARAM = 48842;
      end
      4601: begin
        W_PARAM = 48921;
      end
      4602: begin
        W_PARAM = 16034;
      end
      4603: begin
        W_PARAM = 48484;
      end
      4604: begin
        W_PARAM = 15949;
      end
      4605: begin
        W_PARAM = 15231;
      end
      4606: begin
        W_PARAM = 48726;
      end
      4607: begin
        W_PARAM = 15642;
      end
      4608: begin
        W_PARAM = 16222;
      end
      4609: begin
        W_PARAM = 48682;
      end
      4610: begin
        W_PARAM = 49081;
      end
      4611: begin
        W_PARAM = 16110;
      end
      4612: begin
        W_PARAM = 16169;
      end
      4613: begin
        W_PARAM = 16192;
      end
      4614: begin
        W_PARAM = 48686;
      end
      4615: begin
        W_PARAM = 48661;
      end
      4616: begin
        W_PARAM = 48622;
      end
      4617: begin
        W_PARAM = 15904;
      end
      4618: begin
        W_PARAM = 15798;
      end
      4619: begin
        W_PARAM = 48760;
      end
      4620: begin
        W_PARAM = 48906;
      end
      4621: begin
        W_PARAM = 16240;
      end
      4622: begin
        W_PARAM = 16008;
      end
      4623: begin
        W_PARAM = 15176;
      end
      4624: begin
        W_PARAM = 16137;
      end
      4625: begin
        W_PARAM = 48911;
      end
      4626: begin
        W_PARAM = 15878;
      end
      4627: begin
        W_PARAM = 49015;
      end
      4628: begin
        W_PARAM = 15838;
      end
      4629: begin
        W_PARAM = 15782;
      end
      4630: begin
        W_PARAM = 48696;
      end
      4631: begin
        W_PARAM = 48900;
      end
      4632: begin
        W_PARAM = 48807;
      end
      4633: begin
        W_PARAM = 48624;
      end
      4634: begin
        W_PARAM = 16180;
      end
      4635: begin
        W_PARAM = 48454;
      end
      4636: begin
        W_PARAM = 15857;
      end
      4637: begin
        W_PARAM = 16037;
      end
      4638: begin
        W_PARAM = 15549;
      end
      4639: begin
        W_PARAM = 15505;
      end
      4640: begin
        W_PARAM = 48874;
      end
      4641: begin
        W_PARAM = 16062;
      end
      4642: begin
        W_PARAM = 15917;
      end
      4643: begin
        W_PARAM = 48959;
      end
      4644: begin
        W_PARAM = 16129;
      end
      4645: begin
        W_PARAM = 48844;
      end
      4646: begin
        W_PARAM = 15868;
      end
      4647: begin
        W_PARAM = 48171;
      end
      4648: begin
        W_PARAM = 15984;
      end
      4649: begin
        W_PARAM = 15963;
      end
      4650: begin
        W_PARAM = 15916;
      end
      4651: begin
        W_PARAM = 49101;
      end
      4652: begin
        W_PARAM = 16236;
      end
      4653: begin
        W_PARAM = 48663;
      end
      4654: begin
        W_PARAM = 16065;
      end
      4655: begin
        W_PARAM = 48654;
      end
      4656: begin
        W_PARAM = 48889;
      end
      4657: begin
        W_PARAM = 16112;
      end
      4658: begin
        W_PARAM = 15885;
      end
      4659: begin
        W_PARAM = 16024;
      end
      4660: begin
        W_PARAM = 48163;
      end
      4661: begin
        W_PARAM = 48994;
      end
      4662: begin
        W_PARAM = 48270;
      end
      4663: begin
        W_PARAM = 16169;
      end
      4664: begin
        W_PARAM = 15833;
      end
      4665: begin
        W_PARAM = 48876;
      end
      4666: begin
        W_PARAM = 15910;
      end
      4667: begin
        W_PARAM = 15868;
      end
      4668: begin
        W_PARAM = 15254;
      end
      4669: begin
        W_PARAM = 16034;
      end
      4670: begin
        W_PARAM = 15410;
      end
      4671: begin
        W_PARAM = 48962;
      end
      4672: begin
        W_PARAM = 15531;
      end
      4673: begin
        W_PARAM = 16131;
      end
      4674: begin
        W_PARAM = 15910;
      end
      4675: begin
        W_PARAM = 15861;
      end
      4676: begin
        W_PARAM = 16090;
      end
      4677: begin
        W_PARAM = 16169;
      end
      4678: begin
        W_PARAM = 49003;
      end
      4679: begin
        W_PARAM = 48758;
      end
      4680: begin
        W_PARAM = 16044;
      end
      4681: begin
        W_PARAM = 48797;
      end
      4682: begin
        W_PARAM = 48815;
      end
      4683: begin
        W_PARAM = 15949;
      end
      4684: begin
        W_PARAM = 16186;
      end
      4685: begin
        W_PARAM = 16044;
      end
      4686: begin
        W_PARAM = 48793;
      end
      4687: begin
        W_PARAM = 16008;
      end
      4688: begin
        W_PARAM = 48997;
      end
      4689: begin
        W_PARAM = 48288;
      end
      4690: begin
        W_PARAM = 16001;
      end
      4691: begin
        W_PARAM = 48666;
      end
      4692: begin
        W_PARAM = 16229;
      end
      4693: begin
        W_PARAM = 48556;
      end
      4694: begin
        W_PARAM = 16055;
      end
      4695: begin
        W_PARAM = 48730;
      end
      4696: begin
        W_PARAM = 15957;
      end
      4697: begin
        W_PARAM = 16119;
      end
      4698: begin
        W_PARAM = 49027;
      end
      4699: begin
        W_PARAM = 48953;
      end
      4700: begin
        W_PARAM = 15942;
      end
      4701: begin
        W_PARAM = 48816;
      end
      4702: begin
        W_PARAM = 16133;
      end
      4703: begin
        W_PARAM = 15754;
      end
      4704: begin
        W_PARAM = 48785;
      end
      4705: begin
        W_PARAM = 16180;
      end
      4706: begin
        W_PARAM = 48686;
      end
      4707: begin
        W_PARAM = 48854;
      end
      4708: begin
        W_PARAM = 48933;
      end
      4709: begin
        W_PARAM = 16065;
      end
      4710: begin
        W_PARAM = 48596;
      end
      4711: begin
        W_PARAM = 48834;
      end
      4712: begin
        W_PARAM = 16190;
      end
      4713: begin
        W_PARAM = 16190;
      end
      4714: begin
        W_PARAM = 48679;
      end
      4715: begin
        W_PARAM = 16006;
      end
      4716: begin
        W_PARAM = 48879;
      end
      4717: begin
        W_PARAM = 48797;
      end
      4718: begin
        W_PARAM = 16096;
      end
      4719: begin
        W_PARAM = 48964;
      end
      4720: begin
        W_PARAM = 15865;
      end
      4721: begin
        W_PARAM = 15745;
      end
      4722: begin
        W_PARAM = 16171;
      end
      4723: begin
        W_PARAM = 16290;
      end
      4724: begin
        W_PARAM = 48942;
      end
      4725: begin
        W_PARAM = 48287;
      end
      4726: begin
        W_PARAM = 16072;
      end
      4727: begin
        W_PARAM = 48863;
      end
      4728: begin
        W_PARAM = 48804;
      end
      4729: begin
        W_PARAM = 49031;
      end
      4730: begin
        W_PARAM = 48738;
      end
      4731: begin
        W_PARAM = 48722;
      end
      4732: begin
        W_PARAM = 16390;
      end
      4733: begin
        W_PARAM = 48858;
      end
      4734: begin
        W_PARAM = 48392;
      end
      4735: begin
        W_PARAM = 48843;
      end
      4736: begin
        W_PARAM = 16151;
      end
      4737: begin
        W_PARAM = 48965;
      end
      4738: begin
        W_PARAM = 48715;
      end
      4739: begin
        W_PARAM = 48864;
      end
      4740: begin
        W_PARAM = 48641;
      end
      4741: begin
        W_PARAM = 48571;
      end
      4742: begin
        W_PARAM = 16343;
      end
      4743: begin
        W_PARAM = 48392;
      end
      4744: begin
        W_PARAM = 48772;
      end
      4745: begin
        W_PARAM = 48812;
      end
      4746: begin
        W_PARAM = 48845;
      end
      4747: begin
        W_PARAM = 48709;
      end
      4748: begin
        W_PARAM = 48692;
      end
      4749: begin
        W_PARAM = 48528;
      end
      4750: begin
        W_PARAM = 15275;
      end
      4751: begin
        W_PARAM = 48168;
      end
      4752: begin
        W_PARAM = 16058;
      end
      4753: begin
        W_PARAM = 47885;
      end
      4754: begin
        W_PARAM = 48282;
      end
      4755: begin
        W_PARAM = 48674;
      end
      4756: begin
        W_PARAM = 48672;
      end
      4757: begin
        W_PARAM = 48256;
      end
      4758: begin
        W_PARAM = 48076;
      end
      4759: begin
        W_PARAM = 47756;
      end
      4760: begin
        W_PARAM = 0;
      end
      4761: begin
        W_PARAM = 0;
      end
      4762: begin
        W_PARAM = 0;
      end
      4763: begin
        W_PARAM = 0;
      end
      4764: begin
        W_PARAM = 0;
      end
      4765: begin
        W_PARAM = 0;
      end
      4766: begin
        W_PARAM = 0;
      end
      4767: begin
        W_PARAM = 0;
      end
      4768: begin
        W_PARAM = 0;
      end
      4769: begin
        W_PARAM = 0;
      end
      4770: begin
        W_PARAM = 47048;
      end
      4771: begin
        W_PARAM = 15028;
      end
      4772: begin
        W_PARAM = 48350;
      end
      4773: begin
        W_PARAM = 15600;
      end
      4774: begin
        W_PARAM = 46565;
      end
      4775: begin
        W_PARAM = 47763;
      end
      4776: begin
        W_PARAM = 46890;
      end
      4777: begin
        W_PARAM = 47323;
      end
      4778: begin
        W_PARAM = 47827;
      end
      4779: begin
        W_PARAM = 47661;
      end
      4780: begin
        W_PARAM = 48571;
      end
      4781: begin
        W_PARAM = 14826;
      end
      4782: begin
        W_PARAM = 15955;
      end
      4783: begin
        W_PARAM = 15917;
      end
      4784: begin
        W_PARAM = 15820;
      end
      4785: begin
        W_PARAM = 48693;
      end
      4786: begin
        W_PARAM = 47982;
      end
      4787: begin
        W_PARAM = 48067;
      end
      4788: begin
        W_PARAM = 48102;
      end
      4789: begin
        W_PARAM = 48707;
      end
      4790: begin
        W_PARAM = 48648;
      end
      4791: begin
        W_PARAM = 48012;
      end
      4792: begin
        W_PARAM = 16197;
      end
      4793: begin
        W_PARAM = 16191;
      end
      4794: begin
        W_PARAM = 48971;
      end
      4795: begin
        W_PARAM = 15958;
      end
      4796: begin
        W_PARAM = 48711;
      end
      4797: begin
        W_PARAM = 48775;
      end
      4798: begin
        W_PARAM = 48530;
      end
      4799: begin
        W_PARAM = 48776;
      end
      4800: begin
        W_PARAM = 16017;
      end
      4801: begin
        W_PARAM = 48370;
      end
      4802: begin
        W_PARAM = 16092;
      end
      4803: begin
        W_PARAM = 16246;
      end
      4804: begin
        W_PARAM = 48784;
      end
      4805: begin
        W_PARAM = 15997;
      end
      4806: begin
        W_PARAM = 49006;
      end
      4807: begin
        W_PARAM = 15752;
      end
      4808: begin
        W_PARAM = 48704;
      end
      4809: begin
        W_PARAM = 48911;
      end
      4810: begin
        W_PARAM = 16127;
      end
      4811: begin
        W_PARAM = 48899;
      end
      4812: begin
        W_PARAM = 16036;
      end
      4813: begin
        W_PARAM = 48294;
      end
      4814: begin
        W_PARAM = 48842;
      end
      4815: begin
        W_PARAM = 16084;
      end
      4816: begin
        W_PARAM = 16014;
      end
      4817: begin
        W_PARAM = 15797;
      end
      4818: begin
        W_PARAM = 48835;
      end
      4819: begin
        W_PARAM = 48790;
      end
      4820: begin
        W_PARAM = 16138;
      end
      4821: begin
        W_PARAM = 48959;
      end
      4822: begin
        W_PARAM = 16086;
      end
      4823: begin
        W_PARAM = 15546;
      end
      4824: begin
        W_PARAM = 48706;
      end
      4825: begin
        W_PARAM = 16240;
      end
      4826: begin
        W_PARAM = 15643;
      end
      4827: begin
        W_PARAM = 48793;
      end
      4828: begin
        W_PARAM = 48641;
      end
      4829: begin
        W_PARAM = 48919;
      end
      4830: begin
        W_PARAM = 16132;
      end
      4831: begin
        W_PARAM = 48856;
      end
      4832: begin
        W_PARAM = 15994;
      end
      4833: begin
        W_PARAM = 15936;
      end
      4834: begin
        W_PARAM = 15885;
      end
      4835: begin
        W_PARAM = 48806;
      end
      4836: begin
        W_PARAM = 48680;
      end
      4837: begin
        W_PARAM = 48909;
      end
      4838: begin
        W_PARAM = 15858;
      end
      4839: begin
        W_PARAM = 16005;
      end
      4840: begin
        W_PARAM = 48783;
      end
      4841: begin
        W_PARAM = 48674;
      end
      4842: begin
        W_PARAM = 15884;
      end
      4843: begin
        W_PARAM = 48804;
      end
      4844: begin
        W_PARAM = 16052;
      end
      4845: begin
        W_PARAM = 48786;
      end
      4846: begin
        W_PARAM = 16124;
      end
      4847: begin
        W_PARAM = 48828;
      end
      4848: begin
        W_PARAM = 15765;
      end
      4849: begin
        W_PARAM = 16055;
      end
      4850: begin
        W_PARAM = 16075;
      end
      4851: begin
        W_PARAM = 48840;
      end
      4852: begin
        W_PARAM = 15892;
      end
      4853: begin
        W_PARAM = 49003;
      end
      4854: begin
        W_PARAM = 15929;
      end
      4855: begin
        W_PARAM = 48705;
      end
      4856: begin
        W_PARAM = 16130;
      end
      4857: begin
        W_PARAM = 48675;
      end
      4858: begin
        W_PARAM = 16168;
      end
      4859: begin
        W_PARAM = 48749;
      end
      4860: begin
        W_PARAM = 16162;
      end
      4861: begin
        W_PARAM = 15939;
      end
      4862: begin
        W_PARAM = 16182;
      end
      4863: begin
        W_PARAM = 48985;
      end
      4864: begin
        W_PARAM = 15918;
      end
      4865: begin
        W_PARAM = 48922;
      end
      4866: begin
        W_PARAM = 16233;
      end
      4867: begin
        W_PARAM = 49042;
      end
      4868: begin
        W_PARAM = 48785;
      end
      4869: begin
        W_PARAM = 16005;
      end
      4870: begin
        W_PARAM = 48215;
      end
      4871: begin
        W_PARAM = 48684;
      end
      4872: begin
        W_PARAM = 16014;
      end
      4873: begin
        W_PARAM = 48901;
      end
      4874: begin
        W_PARAM = 15858;
      end
      4875: begin
        W_PARAM = 48829;
      end
      4876: begin
        W_PARAM = 16232;
      end
      4877: begin
        W_PARAM = 48674;
      end
      4878: begin
        W_PARAM = 16079;
      end
      4879: begin
        W_PARAM = 48884;
      end
      4880: begin
        W_PARAM = 15857;
      end
      4881: begin
        W_PARAM = 16045;
      end
      4882: begin
        W_PARAM = 16073;
      end
      4883: begin
        W_PARAM = 48781;
      end
      4884: begin
        W_PARAM = 48804;
      end
      4885: begin
        W_PARAM = 48968;
      end
      4886: begin
        W_PARAM = 48479;
      end
      4887: begin
        W_PARAM = 15423;
      end
      4888: begin
        W_PARAM = 16023;
      end
      4889: begin
        W_PARAM = 16012;
      end
      4890: begin
        W_PARAM = 49009;
      end
      4891: begin
        W_PARAM = 16181;
      end
      4892: begin
        W_PARAM = 16145;
      end
      4893: begin
        W_PARAM = 48815;
      end
      4894: begin
        W_PARAM = 15868;
      end
      4895: begin
        W_PARAM = 48948;
      end
      4896: begin
        W_PARAM = 15939;
      end
      4897: begin
        W_PARAM = 15323;
      end
      4898: begin
        W_PARAM = 16029;
      end
      4899: begin
        W_PARAM = 15786;
      end
      4900: begin
        W_PARAM = 48928;
      end
      4901: begin
        W_PARAM = 16199;
      end
      4902: begin
        W_PARAM = 48141;
      end
      4903: begin
        W_PARAM = 48888;
      end
      4904: begin
        W_PARAM = 16145;
      end
      4905: begin
        W_PARAM = 48845;
      end
      4906: begin
        W_PARAM = 15997;
      end
      4907: begin
        W_PARAM = 15990;
      end
      4908: begin
        W_PARAM = 15750;
      end
      4909: begin
        W_PARAM = 48833;
      end
      4910: begin
        W_PARAM = 48916;
      end
      4911: begin
        W_PARAM = 15981;
      end
      4912: begin
        W_PARAM = 16065;
      end
      4913: begin
        W_PARAM = 48942;
      end
      4914: begin
        W_PARAM = 16104;
      end
      4915: begin
        W_PARAM = 48559;
      end
      4916: begin
        W_PARAM = 15125;
      end
      4917: begin
        W_PARAM = 15989;
      end
      4918: begin
        W_PARAM = 48875;
      end
      4919: begin
        W_PARAM = 16128;
      end
      4920: begin
        W_PARAM = 48702;
      end
      4921: begin
        W_PARAM = 48770;
      end
      4922: begin
        W_PARAM = 15908;
      end
      4923: begin
        W_PARAM = 15658;
      end
      4924: begin
        W_PARAM = 16029;
      end
      4925: begin
        W_PARAM = 48456;
      end
      4926: begin
        W_PARAM = 48699;
      end
      4927: begin
        W_PARAM = 48788;
      end
      4928: begin
        W_PARAM = 16099;
      end
      4929: begin
        W_PARAM = 15379;
      end
      4930: begin
        W_PARAM = 16107;
      end
      4931: begin
        W_PARAM = 49061;
      end
      4932: begin
        W_PARAM = 48911;
      end
      4933: begin
        W_PARAM = 16143;
      end
      4934: begin
        W_PARAM = 16021;
      end
      4935: begin
        W_PARAM = 16079;
      end
      4936: begin
        W_PARAM = 15961;
      end
      4937: begin
        W_PARAM = 48516;
      end
      4938: begin
        W_PARAM = 48691;
      end
      4939: begin
        W_PARAM = 15907;
      end
      4940: begin
        W_PARAM = 48783;
      end
      4941: begin
        W_PARAM = 48699;
      end
      4942: begin
        W_PARAM = 15746;
      end
      4943: begin
        W_PARAM = 48701;
      end
      4944: begin
        W_PARAM = 16170;
      end
      4945: begin
        W_PARAM = 16139;
      end
      4946: begin
        W_PARAM = 15724;
      end
      4947: begin
        W_PARAM = 16022;
      end
      4948: begin
        W_PARAM = 49000;
      end
      4949: begin
        W_PARAM = 48528;
      end
      4950: begin
        W_PARAM = 15995;
      end
      4951: begin
        W_PARAM = 48613;
      end
      4952: begin
        W_PARAM = 15809;
      end
      4953: begin
        W_PARAM = 16135;
      end
      4954: begin
        W_PARAM = 48912;
      end
      4955: begin
        W_PARAM = 16024;
      end
      4956: begin
        W_PARAM = 15998;
      end
      4957: begin
        W_PARAM = 48921;
      end
      4958: begin
        W_PARAM = 15988;
      end
      4959: begin
        W_PARAM = 48835;
      end
      4960: begin
        W_PARAM = 16139;
      end
      4961: begin
        W_PARAM = 48686;
      end
      4962: begin
        W_PARAM = 48660;
      end
      4963: begin
        W_PARAM = 48671;
      end
      4964: begin
        W_PARAM = 15609;
      end
      4965: begin
        W_PARAM = 15269;
      end
      4966: begin
        W_PARAM = 48264;
      end
      4967: begin
        W_PARAM = 15978;
      end
      4968: begin
        W_PARAM = 48499;
      end
      4969: begin
        W_PARAM = 48773;
      end
      4970: begin
        W_PARAM = 48695;
      end
      4971: begin
        W_PARAM = 48700;
      end
      4972: begin
        W_PARAM = 48805;
      end
      4973: begin
        W_PARAM = 47893;
      end
      4974: begin
        W_PARAM = 15947;
      end
      4975: begin
        W_PARAM = 15719;
      end
      4976: begin
        W_PARAM = 16051;
      end
      4977: begin
        W_PARAM = 48643;
      end
      4978: begin
        W_PARAM = 16060;
      end
      4979: begin
        W_PARAM = 48673;
      end
      4980: begin
        W_PARAM = 16038;
      end
      4981: begin
        W_PARAM = 15900;
      end
      4982: begin
        W_PARAM = 15934;
      end
      4983: begin
        W_PARAM = 15879;
      end
      4984: begin
        W_PARAM = 48719;
      end
      4985: begin
        W_PARAM = 48862;
      end
      4986: begin
        W_PARAM = 15996;
      end
      4987: begin
        W_PARAM = 16020;
      end
      4988: begin
        W_PARAM = 48832;
      end
      4989: begin
        W_PARAM = 48803;
      end
      4990: begin
        W_PARAM = 48591;
      end
      4991: begin
        W_PARAM = 15657;
      end
      4992: begin
        W_PARAM = 48812;
      end
      4993: begin
        W_PARAM = 16180;
      end
      4994: begin
        W_PARAM = 48798;
      end
      4995: begin
        W_PARAM = 16058;
      end
      4996: begin
        W_PARAM = 15820;
      end
      4997: begin
        W_PARAM = 48677;
      end
      4998: begin
        W_PARAM = 16159;
      end
      4999: begin
        W_PARAM = 49004;
      end
      5000: begin
        W_PARAM = 15722;
      end
      5001: begin
        W_PARAM = 15913;
      end
      5002: begin
        W_PARAM = 15916;
      end
      5003: begin
        W_PARAM = 48859;
      end
      5004: begin
        W_PARAM = 48963;
      end
      5005: begin
        W_PARAM = 48278;
      end
      5006: begin
        W_PARAM = 16167;
      end
      5007: begin
        W_PARAM = 16141;
      end
      5008: begin
        W_PARAM = 16167;
      end
      5009: begin
        W_PARAM = 49029;
      end
      5010: begin
        W_PARAM = 15754;
      end
      5011: begin
        W_PARAM = 48788;
      end
      5012: begin
        W_PARAM = 16417;
      end
      5013: begin
        W_PARAM = 48958;
      end
      5014: begin
        W_PARAM = 48937;
      end
      5015: begin
        W_PARAM = 48927;
      end
      5016: begin
        W_PARAM = 16162;
      end
      5017: begin
        W_PARAM = 15878;
      end
      5018: begin
        W_PARAM = 48971;
      end
      5019: begin
        W_PARAM = 48758;
      end
      5020: begin
        W_PARAM = 48427;
      end
      5021: begin
        W_PARAM = 15532;
      end
      5022: begin
        W_PARAM = 16185;
      end
      5023: begin
        W_PARAM = 48451;
      end
      5024: begin
        W_PARAM = 48691;
      end
      5025: begin
        W_PARAM = 48604;
      end
      5026: begin
        W_PARAM = 48757;
      end
      5027: begin
        W_PARAM = 15720;
      end
      5028: begin
        W_PARAM = 48675;
      end
      5029: begin
        W_PARAM = 48362;
      end
      5030: begin
        W_PARAM = 15887;
      end
      5031: begin
        W_PARAM = 48289;
      end
      5032: begin
        W_PARAM = 15891;
      end
      5033: begin
        W_PARAM = 47882;
      end
      5034: begin
        W_PARAM = 48662;
      end
      5035: begin
        W_PARAM = 48324;
      end
      5036: begin
        W_PARAM = 48448;
      end
      5037: begin
        W_PARAM = 48415;
      end
      5038: begin
        W_PARAM = 47829;
      end
      5039: begin
        W_PARAM = 47996;
      end
      5040: begin
        W_PARAM = 47119;
      end
      5041: begin
        W_PARAM = 47171;
      end
      5042: begin
        W_PARAM = 47121;
      end
      5043: begin
        W_PARAM = 47833;
      end
      5044: begin
        W_PARAM = 48372;
      end
      5045: begin
        W_PARAM = 47640;
      end
      5046: begin
        W_PARAM = 46530;
      end
      5047: begin
        W_PARAM = 15576;
      end
      5048: begin
        W_PARAM = 47849;
      end
      5049: begin
        W_PARAM = 15349;
      end
      5050: begin
        W_PARAM = 46751;
      end
      5051: begin
        W_PARAM = 14751;
      end
      5052: begin
        W_PARAM = 47818;
      end
      5053: begin
        W_PARAM = 15146;
      end
      5054: begin
        W_PARAM = 46311;
      end
      5055: begin
        W_PARAM = 47666;
      end
      5056: begin
        W_PARAM = 46637;
      end
      5057: begin
        W_PARAM = 14016;
      end
      5058: begin
        W_PARAM = 47620;
      end
      5059: begin
        W_PARAM = 47404;
      end
      5060: begin
        W_PARAM = 48484;
      end
      5061: begin
        W_PARAM = 47815;
      end
      5062: begin
        W_PARAM = 15626;
      end
      5063: begin
        W_PARAM = 15812;
      end
      5064: begin
        W_PARAM = 15716;
      end
      5065: begin
        W_PARAM = 48586;
      end
      5066: begin
        W_PARAM = 47813;
      end
      5067: begin
        W_PARAM = 15804;
      end
      5068: begin
        W_PARAM = 48250;
      end
      5069: begin
        W_PARAM = 48598;
      end
      5070: begin
        W_PARAM = 48690;
      end
      5071: begin
        W_PARAM = 48102;
      end
      5072: begin
        W_PARAM = 16030;
      end
      5073: begin
        W_PARAM = 16264;
      end
      5074: begin
        W_PARAM = 48803;
      end
      5075: begin
        W_PARAM = 15804;
      end
      5076: begin
        W_PARAM = 48463;
      end
      5077: begin
        W_PARAM = 48434;
      end
      5078: begin
        W_PARAM = 48844;
      end
      5079: begin
        W_PARAM = 48882;
      end
      5080: begin
        W_PARAM = 15971;
      end
      5081: begin
        W_PARAM = 48657;
      end
      5082: begin
        W_PARAM = 16164;
      end
      5083: begin
        W_PARAM = 15764;
      end
      5084: begin
        W_PARAM = 15959;
      end
      5085: begin
        W_PARAM = 16204;
      end
      5086: begin
        W_PARAM = 48886;
      end
      5087: begin
        W_PARAM = 48672;
      end
      5088: begin
        W_PARAM = 48910;
      end
      5089: begin
        W_PARAM = 48924;
      end
      5090: begin
        W_PARAM = 48781;
      end
      5091: begin
        W_PARAM = 48922;
      end
      5092: begin
        W_PARAM = 16307;
      end
      5093: begin
        W_PARAM = 16108;
      end
      5094: begin
        W_PARAM = 48557;
      end
      5095: begin
        W_PARAM = 16015;
      end
      5096: begin
        W_PARAM = 48925;
      end
      5097: begin
        W_PARAM = 15920;
      end
      5098: begin
        W_PARAM = 48466;
      end
      5099: begin
        W_PARAM = 48943;
      end
      5100: begin
        W_PARAM = 48354;
      end
      5101: begin
        W_PARAM = 49077;
      end
      5102: begin
        W_PARAM = 15934;
      end
      5103: begin
        W_PARAM = 16157;
      end
      5104: begin
        W_PARAM = 48581;
      end
      5105: begin
        W_PARAM = 16181;
      end
      5106: begin
        W_PARAM = 15792;
      end
      5107: begin
        W_PARAM = 48920;
      end
      5108: begin
        W_PARAM = 16027;
      end
      5109: begin
        W_PARAM = 15987;
      end
      5110: begin
        W_PARAM = 48609;
      end
      5111: begin
        W_PARAM = 48983;
      end
      5112: begin
        W_PARAM = 16167;
      end
      5113: begin
        W_PARAM = 48831;
      end
      5114: begin
        W_PARAM = 15981;
      end
      5115: begin
        W_PARAM = 16033;
      end
      5116: begin
        W_PARAM = 16131;
      end
      5117: begin
        W_PARAM = 48833;
      end
      5118: begin
        W_PARAM = 48166;
      end
      5119: begin
        W_PARAM = 14940;
      end
      5120: begin
        W_PARAM = 16171;
      end
      5121: begin
        W_PARAM = 48265;
      end
      5122: begin
        W_PARAM = 48513;
      end
      5123: begin
        W_PARAM = 15635;
      end
      5124: begin
        W_PARAM = 15802;
      end
      5125: begin
        W_PARAM = 48328;
      end
      5126: begin
        W_PARAM = 48184;
      end
      5127: begin
        W_PARAM = 48803;
      end
      5128: begin
        W_PARAM = 15269;
      end
      5129: begin
        W_PARAM = 48828;
      end
      5130: begin
        W_PARAM = 16150;
      end
      5131: begin
        W_PARAM = 48304;
      end
      5132: begin
        W_PARAM = 48640;
      end
      5133: begin
        W_PARAM = 48921;
      end
      5134: begin
        W_PARAM = 16107;
      end
      5135: begin
        W_PARAM = 48824;
      end
      5136: begin
        W_PARAM = 16103;
      end
      5137: begin
        W_PARAM = 48808;
      end
      5138: begin
        W_PARAM = 15949;
      end
      5139: begin
        W_PARAM = 48775;
      end
      5140: begin
        W_PARAM = 16107;
      end
      5141: begin
        W_PARAM = 48824;
      end
      5142: begin
        W_PARAM = 16045;
      end
      5143: begin
        W_PARAM = 48905;
      end
      5144: begin
        W_PARAM = 48938;
      end
      5145: begin
        W_PARAM = 48749;
      end
      5146: begin
        W_PARAM = 15963;
      end
      5147: begin
        W_PARAM = 48772;
      end
      5148: begin
        W_PARAM = 16114;
      end
      5149: begin
        W_PARAM = 16144;
      end
      5150: begin
        W_PARAM = 15744;
      end
      5151: begin
        W_PARAM = 48716;
      end
      5152: begin
        W_PARAM = 15901;
      end
      5153: begin
        W_PARAM = 48883;
      end
      5154: begin
        W_PARAM = 48654;
      end
      5155: begin
        W_PARAM = 48659;
      end
      5156: begin
        W_PARAM = 48821;
      end
      5157: begin
        W_PARAM = 16007;
      end
      5158: begin
        W_PARAM = 16070;
      end
      5159: begin
        W_PARAM = 16098;
      end
      5160: begin
        W_PARAM = 48857;
      end
      5161: begin
        W_PARAM = 15515;
      end
      5162: begin
        W_PARAM = 16155;
      end
      5163: begin
        W_PARAM = 48986;
      end
      5164: begin
        W_PARAM = 16046;
      end
      5165: begin
        W_PARAM = 15691;
      end
      5166: begin
        W_PARAM = 16301;
      end
      5167: begin
        W_PARAM = 48950;
      end
      5168: begin
        W_PARAM = 16104;
      end
      5169: begin
        W_PARAM = 48981;
      end
      5170: begin
        W_PARAM = 49001;
      end
      5171: begin
        W_PARAM = 48792;
      end
      5172: begin
        W_PARAM = 16010;
      end
      5173: begin
        W_PARAM = 48802;
      end
      5174: begin
        W_PARAM = 16163;
      end
      5175: begin
        W_PARAM = 48662;
      end
      5176: begin
        W_PARAM = 16198;
      end
      5177: begin
        W_PARAM = 16065;
      end
      5178: begin
        W_PARAM = 48467;
      end
      5179: begin
        W_PARAM = 48808;
      end
      5180: begin
        W_PARAM = 48820;
      end
      5181: begin
        W_PARAM = 16072;
      end
      5182: begin
        W_PARAM = 15935;
      end
      5183: begin
        W_PARAM = 48831;
      end
      5184: begin
        W_PARAM = 15927;
      end
      5185: begin
        W_PARAM = 15993;
      end
      5186: begin
        W_PARAM = 48684;
      end
      5187: begin
        W_PARAM = 48823;
      end
      5188: begin
        W_PARAM = 48722;
      end
      5189: begin
        W_PARAM = 16105;
      end
      5190: begin
        W_PARAM = 48642;
      end
      5191: begin
        W_PARAM = 48907;
      end
      5192: begin
        W_PARAM = 48715;
      end
      5193: begin
        W_PARAM = 16103;
      end
      5194: begin
        W_PARAM = 15895;
      end
      5195: begin
        W_PARAM = 15762;
      end
      5196: begin
        W_PARAM = 15922;
      end
      5197: begin
        W_PARAM = 48716;
      end
      5198: begin
        W_PARAM = 15695;
      end
      5199: begin
        W_PARAM = 15920;
      end
      5200: begin
        W_PARAM = 15878;
      end
      5201: begin
        W_PARAM = 49037;
      end
      5202: begin
        W_PARAM = 15841;
      end
      5203: begin
        W_PARAM = 16147;
      end
      5204: begin
        W_PARAM = 16151;
      end
      5205: begin
        W_PARAM = 48460;
      end
      5206: begin
        W_PARAM = 15971;
      end
      5207: begin
        W_PARAM = 48527;
      end
      5208: begin
        W_PARAM = 48872;
      end
      5209: begin
        W_PARAM = 15692;
      end
      5210: begin
        W_PARAM = 48678;
      end
      5211: begin
        W_PARAM = 15987;
      end
      5212: begin
        W_PARAM = 16137;
      end
      5213: begin
        W_PARAM = 15722;
      end
      5214: begin
        W_PARAM = 48852;
      end
      5215: begin
        W_PARAM = 15927;
      end
      5216: begin
        W_PARAM = 16007;
      end
      5217: begin
        W_PARAM = 48766;
      end
      5218: begin
        W_PARAM = 48831;
      end
      5219: begin
        W_PARAM = 48535;
      end
      5220: begin
        W_PARAM = 48440;
      end
      5221: begin
        W_PARAM = 16163;
      end
      5222: begin
        W_PARAM = 48453;
      end
      5223: begin
        W_PARAM = 15803;
      end
      5224: begin
        W_PARAM = 48678;
      end
      5225: begin
        W_PARAM = 48876;
      end
      5226: begin
        W_PARAM = 16004;
      end
      5227: begin
        W_PARAM = 48446;
      end
      5228: begin
        W_PARAM = 48637;
      end
      5229: begin
        W_PARAM = 48591;
      end
      5230: begin
        W_PARAM = 48757;
      end
      5231: begin
        W_PARAM = 47899;
      end
      5232: begin
        W_PARAM = 16066;
      end
      5233: begin
        W_PARAM = 15879;
      end
      5234: begin
        W_PARAM = 48596;
      end
      5235: begin
        W_PARAM = 16046;
      end
      5236: begin
        W_PARAM = 48515;
      end
      5237: begin
        W_PARAM = 48650;
      end
      5238: begin
        W_PARAM = 48571;
      end
      5239: begin
        W_PARAM = 48733;
      end
      5240: begin
        W_PARAM = 48956;
      end
      5241: begin
        W_PARAM = 16012;
      end
      5242: begin
        W_PARAM = 15681;
      end
      5243: begin
        W_PARAM = 15976;
      end
      5244: begin
        W_PARAM = 15836;
      end
      5245: begin
        W_PARAM = 48667;
      end
      5246: begin
        W_PARAM = 48246;
      end
      5247: begin
        W_PARAM = 48548;
      end
      5248: begin
        W_PARAM = 15938;
      end
      5249: begin
        W_PARAM = 15885;
      end
      5250: begin
        W_PARAM = 48880;
      end
      5251: begin
        W_PARAM = 15646;
      end
      5252: begin
        W_PARAM = 16054;
      end
      5253: begin
        W_PARAM = 16088;
      end
      5254: begin
        W_PARAM = 16050;
      end
      5255: begin
        W_PARAM = 48568;
      end
      5256: begin
        W_PARAM = 48550;
      end
      5257: begin
        W_PARAM = 15771;
      end
      5258: begin
        W_PARAM = 48888;
      end
      5259: begin
        W_PARAM = 48623;
      end
      5260: begin
        W_PARAM = 16124;
      end
      5261: begin
        W_PARAM = 48510;
      end
      5262: begin
        W_PARAM = 15962;
      end
      5263: begin
        W_PARAM = 16176;
      end
      5264: begin
        W_PARAM = 48954;
      end
      5265: begin
        W_PARAM = 16011;
      end
      5266: begin
        W_PARAM = 48722;
      end
      5267: begin
        W_PARAM = 48552;
      end
      5268: begin
        W_PARAM = 48762;
      end
      5269: begin
        W_PARAM = 48816;
      end
      5270: begin
        W_PARAM = 16014;
      end
      5271: begin
        W_PARAM = 15757;
      end
      5272: begin
        W_PARAM = 16259;
      end
      5273: begin
        W_PARAM = 15970;
      end
      5274: begin
        W_PARAM = 48783;
      end
      5275: begin
        W_PARAM = 16133;
      end
      5276: begin
        W_PARAM = 15896;
      end
      5277: begin
        W_PARAM = 49047;
      end
      5278: begin
        W_PARAM = 16005;
      end
      5279: begin
        W_PARAM = 49031;
      end
      5280: begin
        W_PARAM = 48249;
      end
      5281: begin
        W_PARAM = 16081;
      end
      5282: begin
        W_PARAM = 16313;
      end
      5283: begin
        W_PARAM = 48954;
      end
      5284: begin
        W_PARAM = 48913;
      end
      5285: begin
        W_PARAM = 16096;
      end
      5286: begin
        W_PARAM = 16068;
      end
      5287: begin
        W_PARAM = 48912;
      end
      5288: begin
        W_PARAM = 15848;
      end
      5289: begin
        W_PARAM = 49002;
      end
      5290: begin
        W_PARAM = 48020;
      end
      5291: begin
        W_PARAM = 16055;
      end
      5292: begin
        W_PARAM = 16313;
      end
      5293: begin
        W_PARAM = 48840;
      end
      5294: begin
        W_PARAM = 48943;
      end
      5295: begin
        W_PARAM = 48826;
      end
      5296: begin
        W_PARAM = 16112;
      end
      5297: begin
        W_PARAM = 15510;
      end
      5298: begin
        W_PARAM = 48921;
      end
      5299: begin
        W_PARAM = 48767;
      end
      5300: begin
        W_PARAM = 48362;
      end
      5301: begin
        W_PARAM = 15890;
      end
      5302: begin
        W_PARAM = 15740;
      end
      5303: begin
        W_PARAM = 48417;
      end
      5304: begin
        W_PARAM = 48418;
      end
      5305: begin
        W_PARAM = 48554;
      end
      5306: begin
        W_PARAM = 48539;
      end
      5307: begin
        W_PARAM = 15916;
      end
      5308: begin
        W_PARAM = 48578;
      end
      5309: begin
        W_PARAM = 48170;
      end
      5310: begin
        W_PARAM = 48289;
      end
      5311: begin
        W_PARAM = 46851;
      end
      5312: begin
        W_PARAM = 15878;
      end
      5313: begin
        W_PARAM = 47476;
      end
      5314: begin
        W_PARAM = 46936;
      end
      5315: begin
        W_PARAM = 48488;
      end
      5316: begin
        W_PARAM = 48475;
      end
      5317: begin
        W_PARAM = 46955;
      end
      5318: begin
        W_PARAM = 47466;
      end
      5319: begin
        W_PARAM = 47634;
      end
      5320: begin
        W_PARAM = 44797;
      end
      5321: begin
        W_PARAM = 14670;
      end
      5322: begin
        W_PARAM = 47382;
      end
      5323: begin
        W_PARAM = 46875;
      end
      5324: begin
        W_PARAM = 45410;
      end
      5325: begin
        W_PARAM = 45858;
      end
      5326: begin
        W_PARAM = 46145;
      end
      5327: begin
        W_PARAM = 46563;
      end
      5328: begin
        W_PARAM = 47153;
      end
      5329: begin
        W_PARAM = 46140;
      end
      5330: begin
        W_PARAM = 15635;
      end
      5331: begin
        W_PARAM = 14898;
      end
      5332: begin
        W_PARAM = 48141;
      end
      5333: begin
        W_PARAM = 47690;
      end
      5334: begin
        W_PARAM = 48516;
      end
      5335: begin
        W_PARAM = 47870;
      end
      5336: begin
        W_PARAM = 47968;
      end
      5337: begin
        W_PARAM = 15871;
      end
      5338: begin
        W_PARAM = 48028;
      end
      5339: begin
        W_PARAM = 48542;
      end
      5340: begin
        W_PARAM = 15376;
      end
      5341: begin
        W_PARAM = 14990;
      end
      5342: begin
        W_PARAM = 15572;
      end
      5343: begin
        W_PARAM = 48326;
      end
      5344: begin
        W_PARAM = 15717;
      end
      5345: begin
        W_PARAM = 48523;
      end
      5346: begin
        W_PARAM = 48034;
      end
      5347: begin
        W_PARAM = 15829;
      end
      5348: begin
        W_PARAM = 48381;
      end
      5349: begin
        W_PARAM = 48523;
      end
      5350: begin
        W_PARAM = 48597;
      end
      5351: begin
        W_PARAM = 48161;
      end
      5352: begin
        W_PARAM = 48684;
      end
      5353: begin
        W_PARAM = 16266;
      end
      5354: begin
        W_PARAM = 16125;
      end
      5355: begin
        W_PARAM = 15736;
      end
      5356: begin
        W_PARAM = 48625;
      end
      5357: begin
        W_PARAM = 48754;
      end
      5358: begin
        W_PARAM = 48909;
      end
      5359: begin
        W_PARAM = 48868;
      end
      5360: begin
        W_PARAM = 48096;
      end
      5361: begin
        W_PARAM = 48825;
      end
      5362: begin
        W_PARAM = 16017;
      end
      5363: begin
        W_PARAM = 15936;
      end
      5364: begin
        W_PARAM = 48450;
      end
      5365: begin
        W_PARAM = 16209;
      end
      5366: begin
        W_PARAM = 48623;
      end
      5367: begin
        W_PARAM = 15940;
      end
      5368: begin
        W_PARAM = 48822;
      end
      5369: begin
        W_PARAM = 48919;
      end
      5370: begin
        W_PARAM = 48661;
      end
      5371: begin
        W_PARAM = 49065;
      end
      5372: begin
        W_PARAM = 15489;
      end
      5373: begin
        W_PARAM = 16252;
      end
      5374: begin
        W_PARAM = 16037;
      end
      5375: begin
        W_PARAM = 15777;
      end
      5376: begin
        W_PARAM = 48559;
      end
      5377: begin
        W_PARAM = 15664;
      end
      5378: begin
        W_PARAM = 16122;
      end
      5379: begin
        W_PARAM = 48834;
      end
      5380: begin
        W_PARAM = 16094;
      end
      5381: begin
        W_PARAM = 48823;
      end
      5382: begin
        W_PARAM = 48764;
      end
      5383: begin
        W_PARAM = 48825;
      end
      5384: begin
        W_PARAM = 48469;
      end
      5385: begin
        W_PARAM = 16119;
      end
      5386: begin
        W_PARAM = 15853;
      end
      5387: begin
        W_PARAM = 48735;
      end
      5388: begin
        W_PARAM = 15805;
      end
      5389: begin
        W_PARAM = 15842;
      end
      5390: begin
        W_PARAM = 16004;
      end
      5391: begin
        W_PARAM = 16189;
      end
      5392: begin
        W_PARAM = 15950;
      end
      5393: begin
        W_PARAM = 48823;
      end
      5394: begin
        W_PARAM = 48187;
      end
      5395: begin
        W_PARAM = 48530;
      end
      5396: begin
        W_PARAM = 15987;
      end
      5397: begin
        W_PARAM = 48966;
      end
      5398: begin
        W_PARAM = 48866;
      end
      5399: begin
        W_PARAM = 15972;
      end
      5400: begin
        W_PARAM = 15845;
      end
      5401: begin
        W_PARAM = 48545;
      end
      5402: begin
        W_PARAM = 15921;
      end
      5403: begin
        W_PARAM = 48708;
      end
      5404: begin
        W_PARAM = 48802;
      end
      5405: begin
        W_PARAM = 16119;
      end
      5406: begin
        W_PARAM = 48654;
      end
      5407: begin
        W_PARAM = 15403;
      end
      5408: begin
        W_PARAM = 15844;
      end
      5409: begin
        W_PARAM = 48678;
      end
      5410: begin
        W_PARAM = 48676;
      end
      5411: begin
        W_PARAM = 16064;
      end
      5412: begin
        W_PARAM = 16139;
      end
      5413: begin
        W_PARAM = 48088;
      end
      5414: begin
        W_PARAM = 48971;
      end
      5415: begin
        W_PARAM = 15702;
      end
      5416: begin
        W_PARAM = 16133;
      end
      5417: begin
        W_PARAM = 48694;
      end
      5418: begin
        W_PARAM = 16046;
      end
      5419: begin
        W_PARAM = 48945;
      end
      5420: begin
        W_PARAM = 16038;
      end
      5421: begin
        W_PARAM = 48028;
      end
      5422: begin
        W_PARAM = 16161;
      end
      5423: begin
        W_PARAM = 15639;
      end
      5424: begin
        W_PARAM = 48985;
      end
      5425: begin
        W_PARAM = 16064;
      end
      5426: begin
        W_PARAM = 16139;
      end
      5427: begin
        W_PARAM = 49067;
      end
      5428: begin
        W_PARAM = 16129;
      end
      5429: begin
        W_PARAM = 48741;
      end
      5430: begin
        W_PARAM = 16125;
      end
      5431: begin
        W_PARAM = 48872;
      end
      5432: begin
        W_PARAM = 15489;
      end
      5433: begin
        W_PARAM = 48860;
      end
      5434: begin
        W_PARAM = 16100;
      end
      5435: begin
        W_PARAM = 48558;
      end
      5436: begin
        W_PARAM = 16251;
      end
      5437: begin
        W_PARAM = 48646;
      end
      5438: begin
        W_PARAM = 48706;
      end
      5439: begin
        W_PARAM = 48933;
      end
      5440: begin
        W_PARAM = 16135;
      end
      5441: begin
        W_PARAM = 48756;
      end
      5442: begin
        W_PARAM = 48168;
      end
      5443: begin
        W_PARAM = 48742;
      end
      5444: begin
        W_PARAM = 49034;
      end
      5445: begin
        W_PARAM = 15816;
      end
      5446: begin
        W_PARAM = 16160;
      end
      5447: begin
        W_PARAM = 15571;
      end
      5448: begin
        W_PARAM = 15681;
      end
      5449: begin
        W_PARAM = 15981;
      end
      5450: begin
        W_PARAM = 48686;
      end
      5451: begin
        W_PARAM = 16111;
      end
      5452: begin
        W_PARAM = 16182;
      end
      5453: begin
        W_PARAM = 48453;
      end
      5454: begin
        W_PARAM = 48820;
      end
      5455: begin
        W_PARAM = 15873;
      end
      5456: begin
        W_PARAM = 15936;
      end
      5457: begin
        W_PARAM = 48811;
      end
      5458: begin
        W_PARAM = 48778;
      end
      5459: begin
        W_PARAM = 48804;
      end
      5460: begin
        W_PARAM = 48847;
      end
      5461: begin
        W_PARAM = 48883;
      end
      5462: begin
        W_PARAM = 15645;
      end
      5463: begin
        W_PARAM = 48465;
      end
      5464: begin
        W_PARAM = 16187;
      end
      5465: begin
        W_PARAM = 48636;
      end
      5466: begin
        W_PARAM = 16171;
      end
      5467: begin
        W_PARAM = 15982;
      end
      5468: begin
        W_PARAM = 48665;
      end
      5469: begin
        W_PARAM = 48880;
      end
      5470: begin
        W_PARAM = 48743;
      end
      5471: begin
        W_PARAM = 16035;
      end
      5472: begin
        W_PARAM = 16088;
      end
      5473: begin
        W_PARAM = 15469;
      end
      5474: begin
        W_PARAM = 48698;
      end
      5475: begin
        W_PARAM = 15818;
      end
      5476: begin
        W_PARAM = 16060;
      end
      5477: begin
        W_PARAM = 48806;
      end
      5478: begin
        W_PARAM = 48645;
      end
      5479: begin
        W_PARAM = 48824;
      end
      5480: begin
        W_PARAM = 48835;
      end
      5481: begin
        W_PARAM = 16155;
      end
      5482: begin
        W_PARAM = 16067;
      end
      5483: begin
        W_PARAM = 15904;
      end
      5484: begin
        W_PARAM = 48761;
      end
      5485: begin
        W_PARAM = 48686;
      end
      5486: begin
        W_PARAM = 15991;
      end
      5487: begin
        W_PARAM = 48920;
      end
      5488: begin
        W_PARAM = 15846;
      end
      5489: begin
        W_PARAM = 48609;
      end
      5490: begin
        W_PARAM = 15949;
      end
      5491: begin
        W_PARAM = 48819;
      end
      5492: begin
        W_PARAM = 16099;
      end
      5493: begin
        W_PARAM = 16101;
      end
      5494: begin
        W_PARAM = 48800;
      end
      5495: begin
        W_PARAM = 48739;
      end
      5496: begin
        W_PARAM = 16064;
      end
      5497: begin
        W_PARAM = 48851;
      end
      5498: begin
        W_PARAM = 16091;
      end
      5499: begin
        W_PARAM = 48921;
      end
      5500: begin
        W_PARAM = 15748;
      end
      5501: begin
        W_PARAM = 48706;
      end
      5502: begin
        W_PARAM = 16037;
      end
      5503: begin
        W_PARAM = 15999;
      end
      5504: begin
        W_PARAM = 48773;
      end
      5505: begin
        W_PARAM = 15969;
      end
      5506: begin
        W_PARAM = 15802;
      end
      5507: begin
        W_PARAM = 48919;
      end
      5508: begin
        W_PARAM = 15959;
      end
      5509: begin
        W_PARAM = 48622;
      end
      5510: begin
        W_PARAM = 48887;
      end
      5511: begin
        W_PARAM = 15815;
      end
      5512: begin
        W_PARAM = 48777;
      end
      5513: begin
        W_PARAM = 15993;
      end
      5514: begin
        W_PARAM = 48730;
      end
      5515: begin
        W_PARAM = 48762;
      end
      5516: begin
        W_PARAM = 16075;
      end
      5517: begin
        W_PARAM = 16035;
      end
      5518: begin
        W_PARAM = 15507;
      end
      5519: begin
        W_PARAM = 15878;
      end
      5520: begin
        W_PARAM = 15844;
      end
      5521: begin
        W_PARAM = 15599;
      end
      5522: begin
        W_PARAM = 15811;
      end
      5523: begin
        W_PARAM = 48593;
      end
      5524: begin
        W_PARAM = 48859;
      end
      5525: begin
        W_PARAM = 16145;
      end
      5526: begin
        W_PARAM = 48573;
      end
      5527: begin
        W_PARAM = 48597;
      end
      5528: begin
        W_PARAM = 48587;
      end
      5529: begin
        W_PARAM = 15548;
      end
      5530: begin
        W_PARAM = 15906;
      end
      5531: begin
        W_PARAM = 15238;
      end
      5532: begin
        W_PARAM = 15921;
      end
      5533: begin
        W_PARAM = 15986;
      end
      5534: begin
        W_PARAM = 15933;
      end
      5535: begin
        W_PARAM = 16041;
      end
      5536: begin
        W_PARAM = 16040;
      end
      5537: begin
        W_PARAM = 48895;
      end
      5538: begin
        W_PARAM = 48908;
      end
      5539: begin
        W_PARAM = 48828;
      end
      5540: begin
        W_PARAM = 16209;
      end
      5541: begin
        W_PARAM = 15874;
      end
      5542: begin
        W_PARAM = 16158;
      end
      5543: begin
        W_PARAM = 48398;
      end
      5544: begin
        W_PARAM = 49064;
      end
      5545: begin
        W_PARAM = 47988;
      end
      5546: begin
        W_PARAM = 16160;
      end
      5547: begin
        W_PARAM = 48969;
      end
      5548: begin
        W_PARAM = 16156;
      end
      5549: begin
        W_PARAM = 48938;
      end
      5550: begin
        W_PARAM = 15662;
      end
      5551: begin
        W_PARAM = 15875;
      end
      5552: begin
        W_PARAM = 16129;
      end
      5553: begin
        W_PARAM = 16149;
      end
      5554: begin
        W_PARAM = 48978;
      end
      5555: begin
        W_PARAM = 16134;
      end
      5556: begin
        W_PARAM = 16023;
      end
      5557: begin
        W_PARAM = 49069;
      end
      5558: begin
        W_PARAM = 16113;
      end
      5559: begin
        W_PARAM = 48832;
      end
      5560: begin
        W_PARAM = 16043;
      end
      5561: begin
        W_PARAM = 16069;
      end
      5562: begin
        W_PARAM = 16053;
      end
      5563: begin
        W_PARAM = 48716;
      end
      5564: begin
        W_PARAM = 48944;
      end
      5565: begin
        W_PARAM = 16173;
      end
      5566: begin
        W_PARAM = 15715;
      end
      5567: begin
        W_PARAM = 48767;
      end
      5568: begin
        W_PARAM = 48792;
      end
      5569: begin
        W_PARAM = 48830;
      end
      5570: begin
        W_PARAM = 48612;
      end
      5571: begin
        W_PARAM = 16109;
      end
      5572: begin
        W_PARAM = 16324;
      end
      5573: begin
        W_PARAM = 48695;
      end
      5574: begin
        W_PARAM = 48855;
      end
      5575: begin
        W_PARAM = 15620;
      end
      5576: begin
        W_PARAM = 48796;
      end
      5577: begin
        W_PARAM = 48652;
      end
      5578: begin
        W_PARAM = 48945;
      end
      5579: begin
        W_PARAM = 48697;
      end
      5580: begin
        W_PARAM = 48353;
      end
      5581: begin
        W_PARAM = 15891;
      end
      5582: begin
        W_PARAM = 16118;
      end
      5583: begin
        W_PARAM = 48271;
      end
      5584: begin
        W_PARAM = 47844;
      end
      5585: begin
        W_PARAM = 48731;
      end
      5586: begin
        W_PARAM = 48722;
      end
      5587: begin
        W_PARAM = 47909;
      end
      5588: begin
        W_PARAM = 48613;
      end
      5589: begin
        W_PARAM = 48439;
      end
      5590: begin
        W_PARAM = 48028;
      end
      5591: begin
        W_PARAM = 14637;
      end
      5592: begin
        W_PARAM = 15717;
      end
      5593: begin
        W_PARAM = 47341;
      end
      5594: begin
        W_PARAM = 46001;
      end
      5595: begin
        W_PARAM = 48273;
      end
      5596: begin
        W_PARAM = 48393;
      end
      5597: begin
        W_PARAM = 46295;
      end
      5598: begin
        W_PARAM = 47238;
      end
      5599: begin
        W_PARAM = 46097;
      end
      5600: begin
        W_PARAM = 0;
      end
      5601: begin
        W_PARAM = 0;
      end
      5602: begin
        W_PARAM = 0;
      end
      5603: begin
        W_PARAM = 0;
      end
      5604: begin
        W_PARAM = 0;
      end
      5605: begin
        W_PARAM = 0;
      end
      5606: begin
        W_PARAM = 0;
      end
      5607: begin
        W_PARAM = 0;
      end
      5608: begin
        W_PARAM = 0;
      end
      5609: begin
        W_PARAM = 0;
      end
      5610: begin
        W_PARAM = 15803;
      end
      5611: begin
        W_PARAM = 47181;
      end
      5612: begin
        W_PARAM = 48283;
      end
      5613: begin
        W_PARAM = 15261;
      end
      5614: begin
        W_PARAM = 47544;
      end
      5615: begin
        W_PARAM = 48126;
      end
      5616: begin
        W_PARAM = 48122;
      end
      5617: begin
        W_PARAM = 47786;
      end
      5618: begin
        W_PARAM = 48171;
      end
      5619: begin
        W_PARAM = 48459;
      end
      5620: begin
        W_PARAM = 48314;
      end
      5621: begin
        W_PARAM = 48164;
      end
      5622: begin
        W_PARAM = 15946;
      end
      5623: begin
        W_PARAM = 48456;
      end
      5624: begin
        W_PARAM = 15746;
      end
      5625: begin
        W_PARAM = 48339;
      end
      5626: begin
        W_PARAM = 48069;
      end
      5627: begin
        W_PARAM = 48305;
      end
      5628: begin
        W_PARAM = 48465;
      end
      5629: begin
        W_PARAM = 48537;
      end
      5630: begin
        W_PARAM = 48654;
      end
      5631: begin
        W_PARAM = 48414;
      end
      5632: begin
        W_PARAM = 16056;
      end
      5633: begin
        W_PARAM = 16196;
      end
      5634: begin
        W_PARAM = 15961;
      end
      5635: begin
        W_PARAM = 15976;
      end
      5636: begin
        W_PARAM = 48632;
      end
      5637: begin
        W_PARAM = 48816;
      end
      5638: begin
        W_PARAM = 48873;
      end
      5639: begin
        W_PARAM = 48879;
      end
      5640: begin
        W_PARAM = 16088;
      end
      5641: begin
        W_PARAM = 48598;
      end
      5642: begin
        W_PARAM = 16092;
      end
      5643: begin
        W_PARAM = 16244;
      end
      5644: begin
        W_PARAM = 15747;
      end
      5645: begin
        W_PARAM = 48773;
      end
      5646: begin
        W_PARAM = 48766;
      end
      5647: begin
        W_PARAM = 48935;
      end
      5648: begin
        W_PARAM = 48799;
      end
      5649: begin
        W_PARAM = 48792;
      end
      5650: begin
        W_PARAM = 16130;
      end
      5651: begin
        W_PARAM = 49065;
      end
      5652: begin
        W_PARAM = 16168;
      end
      5653: begin
        W_PARAM = 16038;
      end
      5654: begin
        W_PARAM = 48912;
      end
      5655: begin
        W_PARAM = 16187;
      end
      5656: begin
        W_PARAM = 48726;
      end
      5657: begin
        W_PARAM = 48900;
      end
      5658: begin
        W_PARAM = 48710;
      end
      5659: begin
        W_PARAM = 16150;
      end
      5660: begin
        W_PARAM = 16034;
      end
      5661: begin
        W_PARAM = 48703;
      end
      5662: begin
        W_PARAM = 16163;
      end
      5663: begin
        W_PARAM = 16193;
      end
      5664: begin
        W_PARAM = 48758;
      end
      5665: begin
        W_PARAM = 16082;
      end
      5666: begin
        W_PARAM = 48804;
      end
      5667: begin
        W_PARAM = 48965;
      end
      5668: begin
        W_PARAM = 48734;
      end
      5669: begin
        W_PARAM = 48838;
      end
      5670: begin
        W_PARAM = 16010;
      end
      5671: begin
        W_PARAM = 15845;
      end
      5672: begin
        W_PARAM = 16259;
      end
      5673: begin
        W_PARAM = 16081;
      end
      5674: begin
        W_PARAM = 48999;
      end
      5675: begin
        W_PARAM = 48734;
      end
      5676: begin
        W_PARAM = 16184;
      end
      5677: begin
        W_PARAM = 48963;
      end
      5678: begin
        W_PARAM = 16156;
      end
      5679: begin
        W_PARAM = 49057;
      end
      5680: begin
        W_PARAM = 16122;
      end
      5681: begin
        W_PARAM = 16142;
      end
      5682: begin
        W_PARAM = 16035;
      end
      5683: begin
        W_PARAM = 15901;
      end
      5684: begin
        W_PARAM = 49043;
      end
      5685: begin
        W_PARAM = 16094;
      end
      5686: begin
        W_PARAM = 48847;
      end
      5687: begin
        W_PARAM = 48601;
      end
      5688: begin
        W_PARAM = 48389;
      end
      5689: begin
        W_PARAM = 48771;
      end
      5690: begin
        W_PARAM = 16037;
      end
      5691: begin
        W_PARAM = 15909;
      end
      5692: begin
        W_PARAM = 16034;
      end
      5693: begin
        W_PARAM = 16172;
      end
      5694: begin
        W_PARAM = 48803;
      end
      5695: begin
        W_PARAM = 16078;
      end
      5696: begin
        W_PARAM = 16051;
      end
      5697: begin
        W_PARAM = 48952;
      end
      5698: begin
        W_PARAM = 48849;
      end
      5699: begin
        W_PARAM = 48967;
      end
      5700: begin
        W_PARAM = 16098;
      end
      5701: begin
        W_PARAM = 16053;
      end
      5702: begin
        W_PARAM = 16046;
      end
      5703: begin
        W_PARAM = 48719;
      end
      5704: begin
        W_PARAM = 48975;
      end
      5705: begin
        W_PARAM = 15455;
      end
      5706: begin
        W_PARAM = 16240;
      end
      5707: begin
        W_PARAM = 48857;
      end
      5708: begin
        W_PARAM = 16004;
      end
      5709: begin
        W_PARAM = 49000;
      end
      5710: begin
        W_PARAM = 16051;
      end
      5711: begin
        W_PARAM = 16100;
      end
      5712: begin
        W_PARAM = 16193;
      end
      5713: begin
        W_PARAM = 48660;
      end
      5714: begin
        W_PARAM = 48734;
      end
      5715: begin
        W_PARAM = 15951;
      end
      5716: begin
        W_PARAM = 16033;
      end
      5717: begin
        W_PARAM = 48906;
      end
      5718: begin
        W_PARAM = 48746;
      end
      5719: begin
        W_PARAM = 49007;
      end
      5720: begin
        W_PARAM = 16222;
      end
      5721: begin
        W_PARAM = 16068;
      end
      5722: begin
        W_PARAM = 16032;
      end
      5723: begin
        W_PARAM = 48995;
      end
      5724: begin
        W_PARAM = 48793;
      end
      5725: begin
        W_PARAM = 15384;
      end
      5726: begin
        W_PARAM = 16254;
      end
      5727: begin
        W_PARAM = 48732;
      end
      5728: begin
        W_PARAM = 47777;
      end
      5729: begin
        W_PARAM = 49045;
      end
      5730: begin
        W_PARAM = 15975;
      end
      5731: begin
        W_PARAM = 48774;
      end
      5732: begin
        W_PARAM = 15888;
      end
      5733: begin
        W_PARAM = 48546;
      end
      5734: begin
        W_PARAM = 48924;
      end
      5735: begin
        W_PARAM = 15940;
      end
      5736: begin
        W_PARAM = 48674;
      end
      5737: begin
        W_PARAM = 15749;
      end
      5738: begin
        W_PARAM = 16102;
      end
      5739: begin
        W_PARAM = 15631;
      end
      5740: begin
        W_PARAM = 15933;
      end
      5741: begin
        W_PARAM = 15207;
      end
      5742: begin
        W_PARAM = 48788;
      end
      5743: begin
        W_PARAM = 15885;
      end
      5744: begin
        W_PARAM = 48695;
      end
      5745: begin
        W_PARAM = 48711;
      end
      5746: begin
        W_PARAM = 16257;
      end
      5747: begin
        W_PARAM = 15891;
      end
      5748: begin
        W_PARAM = 48938;
      end
      5749: begin
        W_PARAM = 48664;
      end
      5750: begin
        W_PARAM = 15851;
      end
      5751: begin
        W_PARAM = 48778;
      end
      5752: begin
        W_PARAM = 15933;
      end
      5753: begin
        W_PARAM = 48695;
      end
      5754: begin
        W_PARAM = 15770;
      end
      5755: begin
        W_PARAM = 15565;
      end
      5756: begin
        W_PARAM = 16034;
      end
      5757: begin
        W_PARAM = 48878;
      end
      5758: begin
        W_PARAM = 16093;
      end
      5759: begin
        W_PARAM = 48754;
      end
      5760: begin
        W_PARAM = 48841;
      end
      5761: begin
        W_PARAM = 16137;
      end
      5762: begin
        W_PARAM = 48420;
      end
      5763: begin
        W_PARAM = 15888;
      end
      5764: begin
        W_PARAM = 16146;
      end
      5765: begin
        W_PARAM = 16053;
      end
      5766: begin
        W_PARAM = 15658;
      end
      5767: begin
        W_PARAM = 48953;
      end
      5768: begin
        W_PARAM = 48894;
      end
      5769: begin
        W_PARAM = 15385;
      end
      5770: begin
        W_PARAM = 48328;
      end
      5771: begin
        W_PARAM = 16139;
      end
      5772: begin
        W_PARAM = 48822;
      end
      5773: begin
        W_PARAM = 15935;
      end
      5774: begin
        W_PARAM = 15943;
      end
      5775: begin
        W_PARAM = 16077;
      end
      5776: begin
        W_PARAM = 48180;
      end
      5777: begin
        W_PARAM = 49011;
      end
      5778: begin
        W_PARAM = 48047;
      end
      5779: begin
        W_PARAM = 15519;
      end
      5780: begin
        W_PARAM = 15821;
      end
      5781: begin
        W_PARAM = 16163;
      end
      5782: begin
        W_PARAM = 15986;
      end
      5783: begin
        W_PARAM = 16141;
      end
      5784: begin
        W_PARAM = 15883;
      end
      5785: begin
        W_PARAM = 15904;
      end
      5786: begin
        W_PARAM = 16141;
      end
      5787: begin
        W_PARAM = 49113;
      end
      5788: begin
        W_PARAM = 48645;
      end
      5789: begin
        W_PARAM = 48907;
      end
      5790: begin
        W_PARAM = 15927;
      end
      5791: begin
        W_PARAM = 16191;
      end
      5792: begin
        W_PARAM = 16096;
      end
      5793: begin
        W_PARAM = 48228;
      end
      5794: begin
        W_PARAM = 48913;
      end
      5795: begin
        W_PARAM = 16059;
      end
      5796: begin
        W_PARAM = 48815;
      end
      5797: begin
        W_PARAM = 48993;
      end
      5798: begin
        W_PARAM = 15892;
      end
      5799: begin
        W_PARAM = 48527;
      end
      5800: begin
        W_PARAM = 15819;
      end
      5801: begin
        W_PARAM = 16037;
      end
      5802: begin
        W_PARAM = 16142;
      end
      5803: begin
        W_PARAM = 16144;
      end
      5804: begin
        W_PARAM = 48833;
      end
      5805: begin
        W_PARAM = 48673;
      end
      5806: begin
        W_PARAM = 16172;
      end
      5807: begin
        W_PARAM = 49072;
      end
      5808: begin
        W_PARAM = 15993;
      end
      5809: begin
        W_PARAM = 48909;
      end
      5810: begin
        W_PARAM = 15629;
      end
      5811: begin
        W_PARAM = 15614;
      end
      5812: begin
        W_PARAM = 16133;
      end
      5813: begin
        W_PARAM = 15931;
      end
      5814: begin
        W_PARAM = 48684;
      end
      5815: begin
        W_PARAM = 15421;
      end
      5816: begin
        W_PARAM = 15975;
      end
      5817: begin
        W_PARAM = 48973;
      end
      5818: begin
        W_PARAM = 16173;
      end
      5819: begin
        W_PARAM = 48950;
      end
      5820: begin
        W_PARAM = 16076;
      end
      5821: begin
        W_PARAM = 15911;
      end
      5822: begin
        W_PARAM = 16083;
      end
      5823: begin
        W_PARAM = 15917;
      end
      5824: begin
        W_PARAM = 48945;
      end
      5825: begin
        W_PARAM = 16241;
      end
      5826: begin
        W_PARAM = 48848;
      end
      5827: begin
        W_PARAM = 48983;
      end
      5828: begin
        W_PARAM = 16078;
      end
      5829: begin
        W_PARAM = 48908;
      end
      5830: begin
        W_PARAM = 48799;
      end
      5831: begin
        W_PARAM = 15666;
      end
      5832: begin
        W_PARAM = 15924;
      end
      5833: begin
        W_PARAM = 16153;
      end
      5834: begin
        W_PARAM = 48930;
      end
      5835: begin
        W_PARAM = 15522;
      end
      5836: begin
        W_PARAM = 15996;
      end
      5837: begin
        W_PARAM = 48927;
      end
      5838: begin
        W_PARAM = 16092;
      end
      5839: begin
        W_PARAM = 15704;
      end
      5840: begin
        W_PARAM = 15702;
      end
      5841: begin
        W_PARAM = 15728;
      end
      5842: begin
        W_PARAM = 16263;
      end
      5843: begin
        W_PARAM = 48687;
      end
      5844: begin
        W_PARAM = 48862;
      end
      5845: begin
        W_PARAM = 15611;
      end
      5846: begin
        W_PARAM = 48680;
      end
      5847: begin
        W_PARAM = 48533;
      end
      5848: begin
        W_PARAM = 48941;
      end
      5849: begin
        W_PARAM = 16038;
      end
      5850: begin
        W_PARAM = 48635;
      end
      5851: begin
        W_PARAM = 15886;
      end
      5852: begin
        W_PARAM = 16133;
      end
      5853: begin
        W_PARAM = 48584;
      end
      5854: begin
        W_PARAM = 48880;
      end
      5855: begin
        W_PARAM = 16134;
      end
      5856: begin
        W_PARAM = 48545;
      end
      5857: begin
        W_PARAM = 48750;
      end
      5858: begin
        W_PARAM = 48855;
      end
      5859: begin
        W_PARAM = 15988;
      end
      5860: begin
        W_PARAM = 47849;
      end
      5861: begin
        W_PARAM = 15882;
      end
      5862: begin
        W_PARAM = 15732;
      end
      5863: begin
        W_PARAM = 15530;
      end
      5864: begin
        W_PARAM = 47619;
      end
      5865: begin
        W_PARAM = 48313;
      end
      5866: begin
        W_PARAM = 48402;
      end
      5867: begin
        W_PARAM = 47816;
      end
      5868: begin
        W_PARAM = 48631;
      end
      5869: begin
        W_PARAM = 48387;
      end
      5870: begin
        W_PARAM = 46307;
      end
      5871: begin
        W_PARAM = 14891;
      end
      5872: begin
        W_PARAM = 47632;
      end
      5873: begin
        W_PARAM = 47024;
      end
      5874: begin
        W_PARAM = 47264;
      end
      5875: begin
        W_PARAM = 14944;
      end
      5876: begin
        W_PARAM = 46480;
      end
      5877: begin
        W_PARAM = 46549;
      end
      5878: begin
        W_PARAM = 47712;
      end
      5879: begin
        W_PARAM = 46563;
      end
      5880: begin
        W_PARAM = 45020;
      end
      5881: begin
        W_PARAM = 14857;
      end
      5882: begin
        W_PARAM = 47509;
      end
      5883: begin
        W_PARAM = 47267;
      end
      5884: begin
        W_PARAM = 46047;
      end
      5885: begin
        W_PARAM = 46424;
      end
      5886: begin
        W_PARAM = 46353;
      end
      5887: begin
        W_PARAM = 47115;
      end
      5888: begin
        W_PARAM = 47362;
      end
      5889: begin
        W_PARAM = 46678;
      end
      5890: begin
        W_PARAM = 47147;
      end
      5891: begin
        W_PARAM = 14599;
      end
      5892: begin
        W_PARAM = 14706;
      end
      5893: begin
        W_PARAM = 15380;
      end
      5894: begin
        W_PARAM = 46591;
      end
      5895: begin
        W_PARAM = 48057;
      end
      5896: begin
        W_PARAM = 46993;
      end
      5897: begin
        W_PARAM = 47788;
      end
      5898: begin
        W_PARAM = 47413;
      end
      5899: begin
        W_PARAM = 47889;
      end
      5900: begin
        W_PARAM = 48657;
      end
      5901: begin
        W_PARAM = 48253;
      end
      5902: begin
        W_PARAM = 16077;
      end
      5903: begin
        W_PARAM = 15881;
      end
      5904: begin
        W_PARAM = 14674;
      end
      5905: begin
        W_PARAM = 48582;
      end
      5906: begin
        W_PARAM = 48181;
      end
      5907: begin
        W_PARAM = 48687;
      end
      5908: begin
        W_PARAM = 48430;
      end
      5909: begin
        W_PARAM = 48483;
      end
      5910: begin
        W_PARAM = 48429;
      end
      5911: begin
        W_PARAM = 15346;
      end
      5912: begin
        W_PARAM = 16122;
      end
      5913: begin
        W_PARAM = 16158;
      end
      5914: begin
        W_PARAM = 48665;
      end
      5915: begin
        W_PARAM = 15983;
      end
      5916: begin
        W_PARAM = 48621;
      end
      5917: begin
        W_PARAM = 48877;
      end
      5918: begin
        W_PARAM = 48793;
      end
      5919: begin
        W_PARAM = 48781;
      end
      5920: begin
        W_PARAM = 48480;
      end
      5921: begin
        W_PARAM = 16021;
      end
      5922: begin
        W_PARAM = 15954;
      end
      5923: begin
        W_PARAM = 16108;
      end
      5924: begin
        W_PARAM = 48722;
      end
      5925: begin
        W_PARAM = 16165;
      end
      5926: begin
        W_PARAM = 48866;
      end
      5927: begin
        W_PARAM = 48958;
      end
      5928: begin
        W_PARAM = 15858;
      end
      5929: begin
        W_PARAM = 48782;
      end
      5930: begin
        W_PARAM = 16012;
      end
      5931: begin
        W_PARAM = 16244;
      end
      5932: begin
        W_PARAM = 48207;
      end
      5933: begin
        W_PARAM = 48803;
      end
      5934: begin
        W_PARAM = 15683;
      end
      5935: begin
        W_PARAM = 15904;
      end
      5936: begin
        W_PARAM = 48920;
      end
      5937: begin
        W_PARAM = 48920;
      end
      5938: begin
        W_PARAM = 48670;
      end
      5939: begin
        W_PARAM = 15994;
      end
      5940: begin
        W_PARAM = 15898;
      end
      5941: begin
        W_PARAM = 16154;
      end
      5942: begin
        W_PARAM = 15939;
      end
      5943: begin
        W_PARAM = 16077;
      end
      5944: begin
        W_PARAM = 48982;
      end
      5945: begin
        W_PARAM = 15895;
      end
      5946: begin
        W_PARAM = 48928;
      end
      5947: begin
        W_PARAM = 48933;
      end
      5948: begin
        W_PARAM = 16142;
      end
      5949: begin
        W_PARAM = 15736;
      end
      5950: begin
        W_PARAM = 15985;
      end
      5951: begin
        W_PARAM = 16003;
      end
      5952: begin
        W_PARAM = 15946;
      end
      5953: begin
        W_PARAM = 16081;
      end
      5954: begin
        W_PARAM = 48974;
      end
      5955: begin
        W_PARAM = 16176;
      end
      5956: begin
        W_PARAM = 15479;
      end
      5957: begin
        W_PARAM = 49026;
      end
      5958: begin
        W_PARAM = 16133;
      end
      5959: begin
        W_PARAM = 48895;
      end
      5960: begin
        W_PARAM = 48871;
      end
      5961: begin
        W_PARAM = 16014;
      end
      5962: begin
        W_PARAM = 48869;
      end
      5963: begin
        W_PARAM = 16118;
      end
      5964: begin
        W_PARAM = 16181;
      end
      5965: begin
        W_PARAM = 48225;
      end
      5966: begin
        W_PARAM = 16016;
      end
      5967: begin
        W_PARAM = 48690;
      end
      5968: begin
        W_PARAM = 48771;
      end
      5969: begin
        W_PARAM = 48848;
      end
      5970: begin
        W_PARAM = 48511;
      end
      5971: begin
        W_PARAM = 48548;
      end
      5972: begin
        W_PARAM = 16081;
      end
      5973: begin
        W_PARAM = 48950;
      end
      5974: begin
        W_PARAM = 15790;
      end
      5975: begin
        W_PARAM = 15923;
      end
      5976: begin
        W_PARAM = 16058;
      end
      5977: begin
        W_PARAM = 48941;
      end
      5978: begin
        W_PARAM = 16155;
      end
      5979: begin
        W_PARAM = 48602;
      end
      5980: begin
        W_PARAM = 16041;
      end
      5981: begin
        W_PARAM = 16144;
      end
      5982: begin
        W_PARAM = 15904;
      end
      5983: begin
        W_PARAM = 48513;
      end
      5984: begin
        W_PARAM = 48764;
      end
      5985: begin
        W_PARAM = 48394;
      end
      5986: begin
        W_PARAM = 15597;
      end
      5987: begin
        W_PARAM = 15443;
      end
      5988: begin
        W_PARAM = 48898;
      end
      5989: begin
        W_PARAM = 48756;
      end
      5990: begin
        W_PARAM = 16043;
      end
      5991: begin
        W_PARAM = 48740;
      end
      5992: begin
        W_PARAM = 15942;
      end
      5993: begin
        W_PARAM = 48757;
      end
      5994: begin
        W_PARAM = 15835;
      end
      5995: begin
        W_PARAM = 16056;
      end
      5996: begin
        W_PARAM = 16073;
      end
      5997: begin
        W_PARAM = 48856;
      end
      5998: begin
        W_PARAM = 15844;
      end
      5999: begin
        W_PARAM = 48925;
      end
      6000: begin
        W_PARAM = 16123;
      end
      6001: begin
        W_PARAM = 48458;
      end
      6002: begin
        W_PARAM = 48783;
      end
      6003: begin
        W_PARAM = 48559;
      end
      6004: begin
        W_PARAM = 15852;
      end
      6005: begin
        W_PARAM = 15648;
      end
      6006: begin
        W_PARAM = 16236;
      end
      6007: begin
        W_PARAM = 48754;
      end
      6008: begin
        W_PARAM = 48849;
      end
      6009: begin
        W_PARAM = 48897;
      end
      6010: begin
        W_PARAM = 15606;
      end
      6011: begin
        W_PARAM = 48153;
      end
      6012: begin
        W_PARAM = 16104;
      end
      6013: begin
        W_PARAM = 48466;
      end
      6014: begin
        W_PARAM = 48833;
      end
      6015: begin
        W_PARAM = 15859;
      end
      6016: begin
        W_PARAM = 16188;
      end
      6017: begin
        W_PARAM = 48905;
      end
      6018: begin
        W_PARAM = 16033;
      end
      6019: begin
        W_PARAM = 48941;
      end
      6020: begin
        W_PARAM = 48583;
      end
      6021: begin
        W_PARAM = 16142;
      end
      6022: begin
        W_PARAM = 16015;
      end
      6023: begin
        W_PARAM = 48750;
      end
      6024: begin
        W_PARAM = 48839;
      end
      6025: begin
        W_PARAM = 15948;
      end
      6026: begin
        W_PARAM = 16240;
      end
      6027: begin
        W_PARAM = 48942;
      end
      6028: begin
        W_PARAM = 15775;
      end
      6029: begin
        W_PARAM = 48934;
      end
      6030: begin
        W_PARAM = 48354;
      end
      6031: begin
        W_PARAM = 16034;
      end
      6032: begin
        W_PARAM = 48650;
      end
      6033: begin
        W_PARAM = 15875;
      end
      6034: begin
        W_PARAM = 16019;
      end
      6035: begin
        W_PARAM = 15858;
      end
      6036: begin
        W_PARAM = 15910;
      end
      6037: begin
        W_PARAM = 48631;
      end
      6038: begin
        W_PARAM = 48668;
      end
      6039: begin
        W_PARAM = 48915;
      end
      6040: begin
        W_PARAM = 15934;
      end
      6041: begin
        W_PARAM = 48770;
      end
      6042: begin
        W_PARAM = 15973;
      end
      6043: begin
        W_PARAM = 15953;
      end
      6044: begin
        W_PARAM = 48884;
      end
      6045: begin
        W_PARAM = 48665;
      end
      6046: begin
        W_PARAM = 16054;
      end
      6047: begin
        W_PARAM = 16003;
      end
      6048: begin
        W_PARAM = 48665;
      end
      6049: begin
        W_PARAM = 48712;
      end
      6050: begin
        W_PARAM = 48852;
      end
      6051: begin
        W_PARAM = 48622;
      end
      6052: begin
        W_PARAM = 16164;
      end
      6053: begin
        W_PARAM = 48667;
      end
      6054: begin
        W_PARAM = 15718;
      end
      6055: begin
        W_PARAM = 16046;
      end
      6056: begin
        W_PARAM = 16153;
      end
      6057: begin
        W_PARAM = 48837;
      end
      6058: begin
        W_PARAM = 15814;
      end
      6059: begin
        W_PARAM = 48938;
      end
      6060: begin
        W_PARAM = 48787;
      end
      6061: begin
        W_PARAM = 16213;
      end
      6062: begin
        W_PARAM = 16066;
      end
      6063: begin
        W_PARAM = 15870;
      end
      6064: begin
        W_PARAM = 48817;
      end
      6065: begin
        W_PARAM = 15408;
      end
      6066: begin
        W_PARAM = 16111;
      end
      6067: begin
        W_PARAM = 48864;
      end
      6068: begin
        W_PARAM = 48593;
      end
      6069: begin
        W_PARAM = 48931;
      end
      6070: begin
        W_PARAM = 48878;
      end
      6071: begin
        W_PARAM = 15689;
      end
      6072: begin
        W_PARAM = 16209;
      end
      6073: begin
        W_PARAM = 16135;
      end
      6074: begin
        W_PARAM = 15891;
      end
      6075: begin
        W_PARAM = 48609;
      end
      6076: begin
        W_PARAM = 16012;
      end
      6077: begin
        W_PARAM = 48975;
      end
      6078: begin
        W_PARAM = 48559;
      end
      6079: begin
        W_PARAM = 48813;
      end
      6080: begin
        W_PARAM = 48789;
      end
      6081: begin
        W_PARAM = 16227;
      end
      6082: begin
        W_PARAM = 48311;
      end
      6083: begin
        W_PARAM = 48801;
      end
      6084: begin
        W_PARAM = 48543;
      end
      6085: begin
        W_PARAM = 16102;
      end
      6086: begin
        W_PARAM = 15914;
      end
      6087: begin
        W_PARAM = 48930;
      end
      6088: begin
        W_PARAM = 16006;
      end
      6089: begin
        W_PARAM = 48858;
      end
      6090: begin
        W_PARAM = 48688;
      end
      6091: begin
        W_PARAM = 16193;
      end
      6092: begin
        W_PARAM = 16032;
      end
      6093: begin
        W_PARAM = 48793;
      end
      6094: begin
        W_PARAM = 48668;
      end
      6095: begin
        W_PARAM = 16149;
      end
      6096: begin
        W_PARAM = 48694;
      end
      6097: begin
        W_PARAM = 49002;
      end
      6098: begin
        W_PARAM = 48568;
      end
      6099: begin
        W_PARAM = 15909;
      end
      6100: begin
        W_PARAM = 15880;
      end
      6101: begin
        W_PARAM = 48926;
      end
      6102: begin
        W_PARAM = 16164;
      end
      6103: begin
        W_PARAM = 15675;
      end
      6104: begin
        W_PARAM = 48540;
      end
      6105: begin
        W_PARAM = 16184;
      end
      6106: begin
        W_PARAM = 16086;
      end
      6107: begin
        W_PARAM = 49001;
      end
      6108: begin
        W_PARAM = 16103;
      end
      6109: begin
        W_PARAM = 48973;
      end
      6110: begin
        W_PARAM = 15864;
      end
      6111: begin
        W_PARAM = 48820;
      end
      6112: begin
        W_PARAM = 16275;
      end
      6113: begin
        W_PARAM = 48798;
      end
      6114: begin
        W_PARAM = 16006;
      end
      6115: begin
        W_PARAM = 15994;
      end
      6116: begin
        W_PARAM = 48114;
      end
      6117: begin
        W_PARAM = 48966;
      end
      6118: begin
        W_PARAM = 48643;
      end
      6119: begin
        W_PARAM = 48718;
      end
      6120: begin
        W_PARAM = 48718;
      end
      6121: begin
        W_PARAM = 16021;
      end
      6122: begin
        W_PARAM = 16167;
      end
      6123: begin
        W_PARAM = 48859;
      end
      6124: begin
        W_PARAM = 48786;
      end
      6125: begin
        W_PARAM = 16119;
      end
      6126: begin
        W_PARAM = 48299;
      end
      6127: begin
        W_PARAM = 48581;
      end
      6128: begin
        W_PARAM = 48995;
      end
      6129: begin
        W_PARAM = 16121;
      end
      6130: begin
        W_PARAM = 48589;
      end
      6131: begin
        W_PARAM = 15685;
      end
      6132: begin
        W_PARAM = 16076;
      end
      6133: begin
        W_PARAM = 48581;
      end
      6134: begin
        W_PARAM = 48864;
      end
      6135: begin
        W_PARAM = 16170;
      end
      6136: begin
        W_PARAM = 48667;
      end
      6137: begin
        W_PARAM = 48558;
      end
      6138: begin
        W_PARAM = 48764;
      end
      6139: begin
        W_PARAM = 15278;
      end
      6140: begin
        W_PARAM = 15882;
      end
      6141: begin
        W_PARAM = 15423;
      end
      6142: begin
        W_PARAM = 15480;
      end
      6143: begin
        W_PARAM = 14987;
      end
      6144: begin
        W_PARAM = 48112;
      end
      6145: begin
        W_PARAM = 15560;
      end
      6146: begin
        W_PARAM = 48195;
      end
      6147: begin
        W_PARAM = 48234;
      end
      6148: begin
        W_PARAM = 48403;
      end
      6149: begin
        W_PARAM = 48625;
      end
      6150: begin
        W_PARAM = 14228;
      end
      6151: begin
        W_PARAM = 43680;
      end
      6152: begin
        W_PARAM = 46662;
      end
      6153: begin
        W_PARAM = 46006;
      end
      6154: begin
        W_PARAM = 45097;
      end
      6155: begin
        W_PARAM = 46267;
      end
      6156: begin
        W_PARAM = 45857;
      end
      6157: begin
        W_PARAM = 44631;
      end
      6158: begin
        W_PARAM = 46959;
      end
      6159: begin
        W_PARAM = 45655;
      end
      6160: begin
        W_PARAM = 45013;
      end
      6161: begin
        W_PARAM = 14853;
      end
      6162: begin
        W_PARAM = 47504;
      end
      6163: begin
        W_PARAM = 47262;
      end
      6164: begin
        W_PARAM = 46040;
      end
      6165: begin
        W_PARAM = 46417;
      end
      6166: begin
        W_PARAM = 46348;
      end
      6167: begin
        W_PARAM = 47111;
      end
      6168: begin
        W_PARAM = 47357;
      end
      6169: begin
        W_PARAM = 46671;
      end
      6170: begin
        W_PARAM = 46254;
      end
      6171: begin
        W_PARAM = 14632;
      end
      6172: begin
        W_PARAM = 47291;
      end
      6173: begin
        W_PARAM = 14700;
      end
      6174: begin
        W_PARAM = 45840;
      end
      6175: begin
        W_PARAM = 47327;
      end
      6176: begin
        W_PARAM = 46133;
      end
      6177: begin
        W_PARAM = 47262;
      end
      6178: begin
        W_PARAM = 47142;
      end
      6179: begin
        W_PARAM = 47261;
      end
      6180: begin
        W_PARAM = 48296;
      end
      6181: begin
        W_PARAM = 48254;
      end
      6182: begin
        W_PARAM = 16050;
      end
      6183: begin
        W_PARAM = 15876;
      end
      6184: begin
        W_PARAM = 47256;
      end
      6185: begin
        W_PARAM = 48490;
      end
      6186: begin
        W_PARAM = 48028;
      end
      6187: begin
        W_PARAM = 48791;
      end
      6188: begin
        W_PARAM = 48361;
      end
      6189: begin
        W_PARAM = 48478;
      end
      6190: begin
        W_PARAM = 48663;
      end
      6191: begin
        W_PARAM = 48506;
      end
      6192: begin
        W_PARAM = 16135;
      end
      6193: begin
        W_PARAM = 16170;
      end
      6194: begin
        W_PARAM = 48718;
      end
      6195: begin
        W_PARAM = 15798;
      end
      6196: begin
        W_PARAM = 48525;
      end
      6197: begin
        W_PARAM = 48947;
      end
      6198: begin
        W_PARAM = 48453;
      end
      6199: begin
        W_PARAM = 48483;
      end
      6200: begin
        W_PARAM = 48938;
      end
      6201: begin
        W_PARAM = 15950;
      end
      6202: begin
        W_PARAM = 16130;
      end
      6203: begin
        W_PARAM = 16068;
      end
      6204: begin
        W_PARAM = 48811;
      end
      6205: begin
        W_PARAM = 16172;
      end
      6206: begin
        W_PARAM = 48712;
      end
      6207: begin
        W_PARAM = 48952;
      end
      6208: begin
        W_PARAM = 16004;
      end
      6209: begin
        W_PARAM = 48604;
      end
      6210: begin
        W_PARAM = 15700;
      end
      6211: begin
        W_PARAM = 16391;
      end
      6212: begin
        W_PARAM = 16022;
      end
      6213: begin
        W_PARAM = 48735;
      end
      6214: begin
        W_PARAM = 48911;
      end
      6215: begin
        W_PARAM = 48865;
      end
      6216: begin
        W_PARAM = 48841;
      end
      6217: begin
        W_PARAM = 48321;
      end
      6218: begin
        W_PARAM = 15752;
      end
      6219: begin
        W_PARAM = 48995;
      end
      6220: begin
        W_PARAM = 48560;
      end
      6221: begin
        W_PARAM = 16232;
      end
      6222: begin
        W_PARAM = 16195;
      end
      6223: begin
        W_PARAM = 16028;
      end
      6224: begin
        W_PARAM = 48849;
      end
      6225: begin
        W_PARAM = 48858;
      end
      6226: begin
        W_PARAM = 48988;
      end
      6227: begin
        W_PARAM = 48729;
      end
      6228: begin
        W_PARAM = 15921;
      end
      6229: begin
        W_PARAM = 48669;
      end
      6230: begin
        W_PARAM = 48771;
      end
      6231: begin
        W_PARAM = 15780;
      end
      6232: begin
        W_PARAM = 16090;
      end
      6233: begin
        W_PARAM = 15994;
      end
      6234: begin
        W_PARAM = 48918;
      end
      6235: begin
        W_PARAM = 48615;
      end
      6236: begin
        W_PARAM = 48694;
      end
      6237: begin
        W_PARAM = 16060;
      end
      6238: begin
        W_PARAM = 16008;
      end
      6239: begin
        W_PARAM = 48768;
      end
      6240: begin
        W_PARAM = 16083;
      end
      6241: begin
        W_PARAM = 15962;
      end
      6242: begin
        W_PARAM = 16128;
      end
      6243: begin
        W_PARAM = 48816;
      end
      6244: begin
        W_PARAM = 48901;
      end
      6245: begin
        W_PARAM = 48636;
      end
      6246: begin
        W_PARAM = 48709;
      end
      6247: begin
        W_PARAM = 15926;
      end
      6248: begin
        W_PARAM = 48769;
      end
      6249: begin
        W_PARAM = 15873;
      end
      6250: begin
        W_PARAM = 16033;
      end
      6251: begin
        W_PARAM = 16004;
      end
      6252: begin
        W_PARAM = 16139;
      end
      6253: begin
        W_PARAM = 15914;
      end
      6254: begin
        W_PARAM = 48982;
      end
      6255: begin
        W_PARAM = 15710;
      end
      6256: begin
        W_PARAM = 16002;
      end
      6257: begin
        W_PARAM = 48777;
      end
      6258: begin
        W_PARAM = 48641;
      end
      6259: begin
        W_PARAM = 48826;
      end
      6260: begin
        W_PARAM = 15930;
      end
      6261: begin
        W_PARAM = 48660;
      end
      6262: begin
        W_PARAM = 15889;
      end
      6263: begin
        W_PARAM = 48709;
      end
      6264: begin
        W_PARAM = 48836;
      end
      6265: begin
        W_PARAM = 48810;
      end
      6266: begin
        W_PARAM = 16104;
      end
      6267: begin
        W_PARAM = 48351;
      end
      6268: begin
        W_PARAM = 15797;
      end
      6269: begin
        W_PARAM = 15963;
      end
      6270: begin
        W_PARAM = 15806;
      end
      6271: begin
        W_PARAM = 48832;
      end
      6272: begin
        W_PARAM = 15894;
      end
      6273: begin
        W_PARAM = 16031;
      end
      6274: begin
        W_PARAM = 48776;
      end
      6275: begin
        W_PARAM = 16002;
      end
      6276: begin
        W_PARAM = 48557;
      end
      6277: begin
        W_PARAM = 48882;
      end
      6278: begin
        W_PARAM = 16090;
      end
      6279: begin
        W_PARAM = 48376;
      end
      6280: begin
        W_PARAM = 15922;
      end
      6281: begin
        W_PARAM = 49025;
      end
      6282: begin
        W_PARAM = 15982;
      end
      6283: begin
        W_PARAM = 48577;
      end
      6284: begin
        W_PARAM = 48879;
      end
      6285: begin
        W_PARAM = 15924;
      end
      6286: begin
        W_PARAM = 16092;
      end
      6287: begin
        W_PARAM = 16053;
      end
      6288: begin
        W_PARAM = 15881;
      end
      6289: begin
        W_PARAM = 15765;
      end
      6290: begin
        W_PARAM = 16298;
      end
      6291: begin
        W_PARAM = 48917;
      end
      6292: begin
        W_PARAM = 15799;
      end
      6293: begin
        W_PARAM = 48775;
      end
      6294: begin
        W_PARAM = 48776;
      end
      6295: begin
        W_PARAM = 15951;
      end
      6296: begin
        W_PARAM = 16163;
      end
      6297: begin
        W_PARAM = 48951;
      end
      6298: begin
        W_PARAM = 15746;
      end
      6299: begin
        W_PARAM = 48896;
      end
      6300: begin
        W_PARAM = 48698;
      end
      6301: begin
        W_PARAM = 48710;
      end
      6302: begin
        W_PARAM = 48722;
      end
      6303: begin
        W_PARAM = 48722;
      end
      6304: begin
        W_PARAM = 48754;
      end
      6305: begin
        W_PARAM = 16016;
      end
      6306: begin
        W_PARAM = 48780;
      end
      6307: begin
        W_PARAM = 16042;
      end
      6308: begin
        W_PARAM = 16092;
      end
      6309: begin
        W_PARAM = 16002;
      end
      6310: begin
        W_PARAM = 15916;
      end
      6311: begin
        W_PARAM = 15550;
      end
      6312: begin
        W_PARAM = 48673;
      end
      6313: begin
        W_PARAM = 15948;
      end
      6314: begin
        W_PARAM = 48936;
      end
      6315: begin
        W_PARAM = 16000;
      end
      6316: begin
        W_PARAM = 16192;
      end
      6317: begin
        W_PARAM = 48785;
      end
      6318: begin
        W_PARAM = 16043;
      end
      6319: begin
        W_PARAM = 48929;
      end
      6320: begin
        W_PARAM = 15802;
      end
      6321: begin
        W_PARAM = 48400;
      end
      6322: begin
        W_PARAM = 15720;
      end
      6323: begin
        W_PARAM = 15285;
      end
      6324: begin
        W_PARAM = 48707;
      end
      6325: begin
        W_PARAM = 16050;
      end
      6326: begin
        W_PARAM = 15971;
      end
      6327: begin
        W_PARAM = 48534;
      end
      6328: begin
        W_PARAM = 48685;
      end
      6329: begin
        W_PARAM = 48771;
      end
      6330: begin
        W_PARAM = 15978;
      end
      6331: begin
        W_PARAM = 16055;
      end
      6332: begin
        W_PARAM = 48718;
      end
      6333: begin
        W_PARAM = 16115;
      end
      6334: begin
        W_PARAM = 48595;
      end
      6335: begin
        W_PARAM = 48731;
      end
      6336: begin
        W_PARAM = 15762;
      end
      6337: begin
        W_PARAM = 48815;
      end
      6338: begin
        W_PARAM = 15779;
      end
      6339: begin
        W_PARAM = 48819;
      end
      6340: begin
        W_PARAM = 48711;
      end
      6341: begin
        W_PARAM = 16205;
      end
      6342: begin
        W_PARAM = 15850;
      end
      6343: begin
        W_PARAM = 48669;
      end
      6344: begin
        W_PARAM = 48812;
      end
      6345: begin
        W_PARAM = 16103;
      end
      6346: begin
        W_PARAM = 48600;
      end
      6347: begin
        W_PARAM = 48817;
      end
      6348: begin
        W_PARAM = 15691;
      end
      6349: begin
        W_PARAM = 48785;
      end
      6350: begin
        W_PARAM = 15831;
      end
      6351: begin
        W_PARAM = 16029;
      end
      6352: begin
        W_PARAM = 16018;
      end
      6353: begin
        W_PARAM = 16010;
      end
      6354: begin
        W_PARAM = 16077;
      end
      6355: begin
        W_PARAM = 16035;
      end
      6356: begin
        W_PARAM = 48718;
      end
      6357: begin
        W_PARAM = 48329;
      end
      6358: begin
        W_PARAM = 48848;
      end
      6359: begin
        W_PARAM = 49031;
      end
      6360: begin
        W_PARAM = 48720;
      end
      6361: begin
        W_PARAM = 16237;
      end
      6362: begin
        W_PARAM = 16083;
      end
      6363: begin
        W_PARAM = 16095;
      end
      6364: begin
        W_PARAM = 48905;
      end
      6365: begin
        W_PARAM = 15521;
      end
      6366: begin
        W_PARAM = 16079;
      end
      6367: begin
        W_PARAM = 48940;
      end
      6368: begin
        W_PARAM = 48896;
      end
      6369: begin
        W_PARAM = 48786;
      end
      6370: begin
        W_PARAM = 15674;
      end
      6371: begin
        W_PARAM = 15970;
      end
      6372: begin
        W_PARAM = 48648;
      end
      6373: begin
        W_PARAM = 48714;
      end
      6374: begin
        W_PARAM = 16195;
      end
      6375: begin
        W_PARAM = 48525;
      end
      6376: begin
        W_PARAM = 16096;
      end
      6377: begin
        W_PARAM = 49045;
      end
      6378: begin
        W_PARAM = 16096;
      end
      6379: begin
        W_PARAM = 48814;
      end
      6380: begin
        W_PARAM = 16134;
      end
      6381: begin
        W_PARAM = 48900;
      end
      6382: begin
        W_PARAM = 16119;
      end
      6383: begin
        W_PARAM = 16108;
      end
      6384: begin
        W_PARAM = 15821;
      end
      6385: begin
        W_PARAM = 16004;
      end
      6386: begin
        W_PARAM = 48827;
      end
      6387: begin
        W_PARAM = 48966;
      end
      6388: begin
        W_PARAM = 48501;
      end
      6389: begin
        W_PARAM = 48610;
      end
      6390: begin
        W_PARAM = 16032;
      end
      6391: begin
        W_PARAM = 48762;
      end
      6392: begin
        W_PARAM = 15770;
      end
      6393: begin
        W_PARAM = 48227;
      end
      6394: begin
        W_PARAM = 48603;
      end
      6395: begin
        W_PARAM = 16158;
      end
      6396: begin
        W_PARAM = 48898;
      end
      6397: begin
        W_PARAM = 48986;
      end
      6398: begin
        W_PARAM = 15962;
      end
      6399: begin
        W_PARAM = 16129;
      end
      6400: begin
        W_PARAM = 48739;
      end
      6401: begin
        W_PARAM = 15474;
      end
      6402: begin
        W_PARAM = 16129;
      end
      6403: begin
        W_PARAM = 48802;
      end
      6404: begin
        W_PARAM = 48816;
      end
      6405: begin
        W_PARAM = 16146;
      end
      6406: begin
        W_PARAM = 48710;
      end
      6407: begin
        W_PARAM = 48596;
      end
      6408: begin
        W_PARAM = 48812;
      end
      6409: begin
        W_PARAM = 16091;
      end
      6410: begin
        W_PARAM = 48558;
      end
      6411: begin
        W_PARAM = 15309;
      end
      6412: begin
        W_PARAM = 15927;
      end
      6413: begin
        W_PARAM = 48561;
      end
      6414: begin
        W_PARAM = 48792;
      end
      6415: begin
        W_PARAM = 16044;
      end
      6416: begin
        W_PARAM = 48383;
      end
      6417: begin
        W_PARAM = 48504;
      end
      6418: begin
        W_PARAM = 48529;
      end
      6419: begin
        W_PARAM = 15836;
      end
      6420: begin
        W_PARAM = 15462;
      end
      6421: begin
        W_PARAM = 15587;
      end
      6422: begin
        W_PARAM = 48653;
      end
      6423: begin
        W_PARAM = 15158;
      end
      6424: begin
        W_PARAM = 15539;
      end
      6425: begin
        W_PARAM = 15883;
      end
      6426: begin
        W_PARAM = 15017;
      end
      6427: begin
        W_PARAM = 48085;
      end
      6428: begin
        W_PARAM = 48335;
      end
      6429: begin
        W_PARAM = 48395;
      end
      6430: begin
        W_PARAM = 14345;
      end
      6431: begin
        W_PARAM = 43796;
      end
      6432: begin
        W_PARAM = 46775;
      end
      6433: begin
        W_PARAM = 46120;
      end
      6434: begin
        W_PARAM = 45212;
      end
      6435: begin
        W_PARAM = 46380;
      end
      6436: begin
        W_PARAM = 45973;
      end
      6437: begin
        W_PARAM = 44742;
      end
      6438: begin
        W_PARAM = 47069;
      end
      6439: begin
        W_PARAM = 45767;
      end
      6440: begin
        W_PARAM = 0;
      end
      6441: begin
        W_PARAM = 0;
      end
      6442: begin
        W_PARAM = 0;
      end
      6443: begin
        W_PARAM = 0;
      end
      6444: begin
        W_PARAM = 0;
      end
      6445: begin
        W_PARAM = 0;
      end
      6446: begin
        W_PARAM = 0;
      end
      6447: begin
        W_PARAM = 0;
      end
      6448: begin
        W_PARAM = 0;
      end
      6449: begin
        W_PARAM = 0;
      end
      6450: begin
        W_PARAM = 0;
      end
      6451: begin
        W_PARAM = 0;
      end
      6452: begin
        W_PARAM = 0;
      end
      6453: begin
        W_PARAM = 0;
      end
      6454: begin
        W_PARAM = 0;
      end
      6455: begin
        W_PARAM = 0;
      end
      6456: begin
        W_PARAM = 0;
      end
      6457: begin
        W_PARAM = 0;
      end
      6458: begin
        W_PARAM = 0;
      end
      6459: begin
        W_PARAM = 0;
      end
      6460: begin
        W_PARAM = 47522;
      end
      6461: begin
        W_PARAM = 47512;
      end
      6462: begin
        W_PARAM = 15590;
      end
      6463: begin
        W_PARAM = 16013;
      end
      6464: begin
        W_PARAM = 47377;
      end
      6465: begin
        W_PARAM = 47499;
      end
      6466: begin
        W_PARAM = 46632;
      end
      6467: begin
        W_PARAM = 48724;
      end
      6468: begin
        W_PARAM = 48024;
      end
      6469: begin
        W_PARAM = 48571;
      end
      6470: begin
        W_PARAM = 48534;
      end
      6471: begin
        W_PARAM = 48785;
      end
      6472: begin
        W_PARAM = 48584;
      end
      6473: begin
        W_PARAM = 16241;
      end
      6474: begin
        W_PARAM = 48344;
      end
      6475: begin
        W_PARAM = 15982;
      end
      6476: begin
        W_PARAM = 47795;
      end
      6477: begin
        W_PARAM = 48924;
      end
      6478: begin
        W_PARAM = 48631;
      end
      6479: begin
        W_PARAM = 15652;
      end
      6480: begin
        W_PARAM = 48855;
      end
      6481: begin
        W_PARAM = 48911;
      end
      6482: begin
        W_PARAM = 15913;
      end
      6483: begin
        W_PARAM = 16232;
      end
      6484: begin
        W_PARAM = 48740;
      end
      6485: begin
        W_PARAM = 16172;
      end
      6486: begin
        W_PARAM = 48285;
      end
      6487: begin
        W_PARAM = 48659;
      end
      6488: begin
        W_PARAM = 15654;
      end
      6489: begin
        W_PARAM = 48855;
      end
      6490: begin
        W_PARAM = 48775;
      end
      6491: begin
        W_PARAM = 16196;
      end
      6492: begin
        W_PARAM = 48537;
      end
      6493: begin
        W_PARAM = 16183;
      end
      6494: begin
        W_PARAM = 48852;
      end
      6495: begin
        W_PARAM = 16135;
      end
      6496: begin
        W_PARAM = 48607;
      end
      6497: begin
        W_PARAM = 15515;
      end
      6498: begin
        W_PARAM = 48881;
      end
      6499: begin
        W_PARAM = 48946;
      end
      6500: begin
        W_PARAM = 48634;
      end
      6501: begin
        W_PARAM = 16045;
      end
      6502: begin
        W_PARAM = 15866;
      end
      6503: begin
        W_PARAM = 16078;
      end
      6504: begin
        W_PARAM = 48075;
      end
      6505: begin
        W_PARAM = 16000;
      end
      6506: begin
        W_PARAM = 48791;
      end
      6507: begin
        W_PARAM = 15921;
      end
      6508: begin
        W_PARAM = 48859;
      end
      6509: begin
        W_PARAM = 48863;
      end
      6510: begin
        W_PARAM = 16071;
      end
      6511: begin
        W_PARAM = 15894;
      end
      6512: begin
        W_PARAM = 15829;
      end
      6513: begin
        W_PARAM = 16076;
      end
      6514: begin
        W_PARAM = 15767;
      end
      6515: begin
        W_PARAM = 48920;
      end
      6516: begin
        W_PARAM = 48901;
      end
      6517: begin
        W_PARAM = 16181;
      end
      6518: begin
        W_PARAM = 48798;
      end
      6519: begin
        W_PARAM = 48844;
      end
      6520: begin
        W_PARAM = 15958;
      end
      6521: begin
        W_PARAM = 48605;
      end
      6522: begin
        W_PARAM = 15632;
      end
      6523: begin
        W_PARAM = 15760;
      end
      6524: begin
        W_PARAM = 15766;
      end
      6525: begin
        W_PARAM = 16082;
      end
      6526: begin
        W_PARAM = 48799;
      end
      6527: begin
        W_PARAM = 49038;
      end
      6528: begin
        W_PARAM = 16110;
      end
      6529: begin
        W_PARAM = 16006;
      end
      6530: begin
        W_PARAM = 16106;
      end
      6531: begin
        W_PARAM = 15988;
      end
      6532: begin
        W_PARAM = 16062;
      end
      6533: begin
        W_PARAM = 16036;
      end
      6534: begin
        W_PARAM = 48650;
      end
      6535: begin
        W_PARAM = 48541;
      end
      6536: begin
        W_PARAM = 48796;
      end
      6537: begin
        W_PARAM = 48793;
      end
      6538: begin
        W_PARAM = 15849;
      end
      6539: begin
        W_PARAM = 48944;
      end
      6540: begin
        W_PARAM = 16107;
      end
      6541: begin
        W_PARAM = 48725;
      end
      6542: begin
        W_PARAM = 48571;
      end
      6543: begin
        W_PARAM = 15733;
      end
      6544: begin
        W_PARAM = 15529;
      end
      6545: begin
        W_PARAM = 16183;
      end
      6546: begin
        W_PARAM = 48937;
      end
      6547: begin
        W_PARAM = 48745;
      end
      6548: begin
        W_PARAM = 48593;
      end
      6549: begin
        W_PARAM = 15639;
      end
      6550: begin
        W_PARAM = 16123;
      end
      6551: begin
        W_PARAM = 48557;
      end
      6552: begin
        W_PARAM = 16065;
      end
      6553: begin
        W_PARAM = 16135;
      end
      6554: begin
        W_PARAM = 48553;
      end
      6555: begin
        W_PARAM = 48064;
      end
      6556: begin
        W_PARAM = 48792;
      end
      6557: begin
        W_PARAM = 48927;
      end
      6558: begin
        W_PARAM = 15532;
      end
      6559: begin
        W_PARAM = 48806;
      end
      6560: begin
        W_PARAM = 48171;
      end
      6561: begin
        W_PARAM = 16193;
      end
      6562: begin
        W_PARAM = 16042;
      end
      6563: begin
        W_PARAM = 48931;
      end
      6564: begin
        W_PARAM = 48747;
      end
      6565: begin
        W_PARAM = 47889;
      end
      6566: begin
        W_PARAM = 15968;
      end
      6567: begin
        W_PARAM = 48922;
      end
      6568: begin
        W_PARAM = 16024;
      end
      6569: begin
        W_PARAM = 48631;
      end
      6570: begin
        W_PARAM = 15941;
      end
      6571: begin
        W_PARAM = 15818;
      end
      6572: begin
        W_PARAM = 48831;
      end
      6573: begin
        W_PARAM = 16147;
      end
      6574: begin
        W_PARAM = 48699;
      end
      6575: begin
        W_PARAM = 48759;
      end
      6576: begin
        W_PARAM = 48773;
      end
      6577: begin
        W_PARAM = 48887;
      end
      6578: begin
        W_PARAM = 16198;
      end
      6579: begin
        W_PARAM = 48583;
      end
      6580: begin
        W_PARAM = 16033;
      end
      6581: begin
        W_PARAM = 48906;
      end
      6582: begin
        W_PARAM = 48311;
      end
      6583: begin
        W_PARAM = 48816;
      end
      6584: begin
        W_PARAM = 15898;
      end
      6585: begin
        W_PARAM = 16066;
      end
      6586: begin
        W_PARAM = 16023;
      end
      6587: begin
        W_PARAM = 48895;
      end
      6588: begin
        W_PARAM = 15774;
      end
      6589: begin
        W_PARAM = 15935;
      end
      6590: begin
        W_PARAM = 16053;
      end
      6591: begin
        W_PARAM = 16087;
      end
      6592: begin
        W_PARAM = 48802;
      end
      6593: begin
        W_PARAM = 15821;
      end
      6594: begin
        W_PARAM = 48611;
      end
      6595: begin
        W_PARAM = 48772;
      end
      6596: begin
        W_PARAM = 48344;
      end
      6597: begin
        W_PARAM = 48535;
      end
      6598: begin
        W_PARAM = 15968;
      end
      6599: begin
        W_PARAM = 48797;
      end
      6600: begin
        W_PARAM = 48703;
      end
      6601: begin
        W_PARAM = 48435;
      end
      6602: begin
        W_PARAM = 16012;
      end
      6603: begin
        W_PARAM = 48921;
      end
      6604: begin
        W_PARAM = 16058;
      end
      6605: begin
        W_PARAM = 16118;
      end
      6606: begin
        W_PARAM = 48525;
      end
      6607: begin
        W_PARAM = 48915;
      end
      6608: begin
        W_PARAM = 16125;
      end
      6609: begin
        W_PARAM = 48652;
      end
      6610: begin
        W_PARAM = 16060;
      end
      6611: begin
        W_PARAM = 16156;
      end
      6612: begin
        W_PARAM = 48714;
      end
      6613: begin
        W_PARAM = 48046;
      end
      6614: begin
        W_PARAM = 48779;
      end
      6615: begin
        W_PARAM = 15617;
      end
      6616: begin
        W_PARAM = 15682;
      end
      6617: begin
        W_PARAM = 48783;
      end
      6618: begin
        W_PARAM = 48189;
      end
      6619: begin
        W_PARAM = 48790;
      end
      6620: begin
        W_PARAM = 48952;
      end
      6621: begin
        W_PARAM = 48851;
      end
      6622: begin
        W_PARAM = 16110;
      end
      6623: begin
        W_PARAM = 16188;
      end
      6624: begin
        W_PARAM = 16039;
      end
      6625: begin
        W_PARAM = 48924;
      end
      6626: begin
        W_PARAM = 16036;
      end
      6627: begin
        W_PARAM = 48860;
      end
      6628: begin
        W_PARAM = 16103;
      end
      6629: begin
        W_PARAM = 48645;
      end
      6630: begin
        W_PARAM = 48895;
      end
      6631: begin
        W_PARAM = 15820;
      end
      6632: begin
        W_PARAM = 16185;
      end
      6633: begin
        W_PARAM = 48772;
      end
      6634: begin
        W_PARAM = 15874;
      end
      6635: begin
        W_PARAM = 48735;
      end
      6636: begin
        W_PARAM = 16106;
      end
      6637: begin
        W_PARAM = 49005;
      end
      6638: begin
        W_PARAM = 15983;
      end
      6639: begin
        W_PARAM = 16003;
      end
      6640: begin
        W_PARAM = 48925;
      end
      6641: begin
        W_PARAM = 48747;
      end
      6642: begin
        W_PARAM = 16168;
      end
      6643: begin
        W_PARAM = 16031;
      end
      6644: begin
        W_PARAM = 15965;
      end
      6645: begin
        W_PARAM = 16034;
      end
      6646: begin
        W_PARAM = 16035;
      end
      6647: begin
        W_PARAM = 49041;
      end
      6648: begin
        W_PARAM = 15972;
      end
      6649: begin
        W_PARAM = 48523;
      end
      6650: begin
        W_PARAM = 48761;
      end
      6651: begin
        W_PARAM = 48822;
      end
      6652: begin
        W_PARAM = 16214;
      end
      6653: begin
        W_PARAM = 15551;
      end
      6654: begin
        W_PARAM = 16149;
      end
      6655: begin
        W_PARAM = 47792;
      end
      6656: begin
        W_PARAM = 15540;
      end
      6657: begin
        W_PARAM = 49049;
      end
      6658: begin
        W_PARAM = 15818;
      end
      6659: begin
        W_PARAM = 15980;
      end
      6660: begin
        W_PARAM = 48508;
      end
      6661: begin
        W_PARAM = 48721;
      end
      6662: begin
        W_PARAM = 16225;
      end
      6663: begin
        W_PARAM = 48903;
      end
      6664: begin
        W_PARAM = 48921;
      end
      6665: begin
        W_PARAM = 15534;
      end
      6666: begin
        W_PARAM = 48452;
      end
      6667: begin
        W_PARAM = 48916;
      end
      6668: begin
        W_PARAM = 15991;
      end
      6669: begin
        W_PARAM = 16224;
      end
      6670: begin
        W_PARAM = 48734;
      end
      6671: begin
        W_PARAM = 48786;
      end
      6672: begin
        W_PARAM = 16169;
      end
      6673: begin
        W_PARAM = 48697;
      end
      6674: begin
        W_PARAM = 48875;
      end
      6675: begin
        W_PARAM = 16062;
      end
      6676: begin
        W_PARAM = 48645;
      end
      6677: begin
        W_PARAM = 48993;
      end
      6678: begin
        W_PARAM = 16115;
      end
      6679: begin
        W_PARAM = 16164;
      end
      6680: begin
        W_PARAM = 48819;
      end
      6681: begin
        W_PARAM = 48551;
      end
      6682: begin
        W_PARAM = 16181;
      end
      6683: begin
        W_PARAM = 48549;
      end
      6684: begin
        W_PARAM = 48821;
      end
      6685: begin
        W_PARAM = 16023;
      end
      6686: begin
        W_PARAM = 48612;
      end
      6687: begin
        W_PARAM = 48769;
      end
      6688: begin
        W_PARAM = 48738;
      end
      6689: begin
        W_PARAM = 16101;
      end
      6690: begin
        W_PARAM = 48488;
      end
      6691: begin
        W_PARAM = 15077;
      end
      6692: begin
        W_PARAM = 16002;
      end
      6693: begin
        W_PARAM = 48578;
      end
      6694: begin
        W_PARAM = 15421;
      end
      6695: begin
        W_PARAM = 15841;
      end
      6696: begin
        W_PARAM = 48272;
      end
      6697: begin
        W_PARAM = 48532;
      end
      6698: begin
        W_PARAM = 48542;
      end
      6699: begin
        W_PARAM = 48491;
      end
      6700: begin
        W_PARAM = 46988;
      end
      6701: begin
        W_PARAM = 15867;
      end
      6702: begin
        W_PARAM = 48569;
      end
      6703: begin
        W_PARAM = 15721;
      end
      6704: begin
        W_PARAM = 15544;
      end
      6705: begin
        W_PARAM = 15782;
      end
      6706: begin
        W_PARAM = 47445;
      end
      6707: begin
        W_PARAM = 48038;
      end
      6708: begin
        W_PARAM = 48619;
      end
      6709: begin
        W_PARAM = 48533;
      end
      6710: begin
        W_PARAM = 0;
      end
      6711: begin
        W_PARAM = 0;
      end
      6712: begin
        W_PARAM = 0;
      end
      6713: begin
        W_PARAM = 0;
      end
      6714: begin
        W_PARAM = 0;
      end
      6715: begin
        W_PARAM = 0;
      end
      6716: begin
        W_PARAM = 0;
      end
      6717: begin
        W_PARAM = 0;
      end
      6718: begin
        W_PARAM = 0;
      end
      6719: begin
        W_PARAM = 0;
      end
      6720: begin
        W_PARAM = 0;
      end
      6721: begin
        W_PARAM = 0;
      end
      6722: begin
        W_PARAM = 0;
      end
      6723: begin
        W_PARAM = 0;
      end
      6724: begin
        W_PARAM = 0;
      end
      6725: begin
        W_PARAM = 0;
      end
      6726: begin
        W_PARAM = 0;
      end
      6727: begin
        W_PARAM = 0;
      end
      6728: begin
        W_PARAM = 0;
      end
      6729: begin
        W_PARAM = 0;
      end
      6730: begin
        W_PARAM = 0;
      end
      6731: begin
        W_PARAM = 0;
      end
      6732: begin
        W_PARAM = 0;
      end
      6733: begin
        W_PARAM = 0;
      end
      6734: begin
        W_PARAM = 0;
      end
      6735: begin
        W_PARAM = 0;
      end
      6736: begin
        W_PARAM = 0;
      end
      6737: begin
        W_PARAM = 0;
      end
      6738: begin
        W_PARAM = 0;
      end
      6739: begin
        W_PARAM = 0;
      end
      6740: begin
        W_PARAM = 47814;
      end
      6741: begin
        W_PARAM = 46636;
      end
      6742: begin
        W_PARAM = 47903;
      end
      6743: begin
        W_PARAM = 15849;
      end
      6744: begin
        W_PARAM = 46903;
      end
      6745: begin
        W_PARAM = 47647;
      end
      6746: begin
        W_PARAM = 46217;
      end
      6747: begin
        W_PARAM = 48564;
      end
      6748: begin
        W_PARAM = 47480;
      end
      6749: begin
        W_PARAM = 48299;
      end
      6750: begin
        W_PARAM = 47889;
      end
      6751: begin
        W_PARAM = 48693;
      end
      6752: begin
        W_PARAM = 48800;
      end
      6753: begin
        W_PARAM = 16142;
      end
      6754: begin
        W_PARAM = 47444;
      end
      6755: begin
        W_PARAM = 16009;
      end
      6756: begin
        W_PARAM = 47089;
      end
      6757: begin
        W_PARAM = 48407;
      end
      6758: begin
        W_PARAM = 48769;
      end
      6759: begin
        W_PARAM = 48425;
      end
      6760: begin
        W_PARAM = 15822;
      end
      6761: begin
        W_PARAM = 48788;
      end
      6762: begin
        W_PARAM = 48865;
      end
      6763: begin
        W_PARAM = 16207;
      end
      6764: begin
        W_PARAM = 48533;
      end
      6765: begin
        W_PARAM = 15300;
      end
      6766: begin
        W_PARAM = 47915;
      end
      6767: begin
        W_PARAM = 16002;
      end
      6768: begin
        W_PARAM = 48921;
      end
      6769: begin
        W_PARAM = 15982;
      end
      6770: begin
        W_PARAM = 48665;
      end
      6771: begin
        W_PARAM = 15570;
      end
      6772: begin
        W_PARAM = 48920;
      end
      6773: begin
        W_PARAM = 15942;
      end
      6774: begin
        W_PARAM = 48356;
      end
      6775: begin
        W_PARAM = 15704;
      end
      6776: begin
        W_PARAM = 48470;
      end
      6777: begin
        W_PARAM = 16258;
      end
      6778: begin
        W_PARAM = 48970;
      end
      6779: begin
        W_PARAM = 16039;
      end
      6780: begin
        W_PARAM = 48825;
      end
      6781: begin
        W_PARAM = 48642;
      end
      6782: begin
        W_PARAM = 48928;
      end
      6783: begin
        W_PARAM = 16219;
      end
      6784: begin
        W_PARAM = 15819;
      end
      6785: begin
        W_PARAM = 48434;
      end
      6786: begin
        W_PARAM = 48534;
      end
      6787: begin
        W_PARAM = 16201;
      end
      6788: begin
        W_PARAM = 48929;
      end
      6789: begin
        W_PARAM = 15863;
      end
      6790: begin
        W_PARAM = 48862;
      end
      6791: begin
        W_PARAM = 48662;
      end
      6792: begin
        W_PARAM = 48883;
      end
      6793: begin
        W_PARAM = 16149;
      end
      6794: begin
        W_PARAM = 15941;
      end
      6795: begin
        W_PARAM = 15856;
      end
      6796: begin
        W_PARAM = 48751;
      end
      6797: begin
        W_PARAM = 16089;
      end
      6798: begin
        W_PARAM = 48773;
      end
      6799: begin
        W_PARAM = 15981;
      end
      6800: begin
        W_PARAM = 48321;
      end
      6801: begin
        W_PARAM = 48825;
      end
      6802: begin
        W_PARAM = 48535;
      end
      6803: begin
        W_PARAM = 48467;
      end
      6804: begin
        W_PARAM = 15427;
      end
      6805: begin
        W_PARAM = 15964;
      end
      6806: begin
        W_PARAM = 48870;
      end
      6807: begin
        W_PARAM = 16009;
      end
      6808: begin
        W_PARAM = 16075;
      end
      6809: begin
        W_PARAM = 15756;
      end
      6810: begin
        W_PARAM = 16029;
      end
      6811: begin
        W_PARAM = 48700;
      end
      6812: begin
        W_PARAM = 16018;
      end
      6813: begin
        W_PARAM = 15881;
      end
      6814: begin
        W_PARAM = 16004;
      end
      6815: begin
        W_PARAM = 16130;
      end
      6816: begin
        W_PARAM = 48929;
      end
      6817: begin
        W_PARAM = 48715;
      end
      6818: begin
        W_PARAM = 48514;
      end
      6819: begin
        W_PARAM = 48855;
      end
      6820: begin
        W_PARAM = 15825;
      end
      6821: begin
        W_PARAM = 48721;
      end
      6822: begin
        W_PARAM = 48517;
      end
      6823: begin
        W_PARAM = 16144;
      end
      6824: begin
        W_PARAM = 48049;
      end
      6825: begin
        W_PARAM = 15750;
      end
      6826: begin
        W_PARAM = 48969;
      end
      6827: begin
        W_PARAM = 15796;
      end
      6828: begin
        W_PARAM = 15642;
      end
      6829: begin
        W_PARAM = 15954;
      end
      6830: begin
        W_PARAM = 48867;
      end
      6831: begin
        W_PARAM = 48686;
      end
      6832: begin
        W_PARAM = 48432;
      end
      6833: begin
        W_PARAM = 16138;
      end
      6834: begin
        W_PARAM = 16167;
      end
      6835: begin
        W_PARAM = 16021;
      end
      6836: begin
        W_PARAM = 49055;
      end
      6837: begin
        W_PARAM = 48669;
      end
      6838: begin
        W_PARAM = 16172;
      end
      6839: begin
        W_PARAM = 48605;
      end
      6840: begin
        W_PARAM = 16188;
      end
      6841: begin
        W_PARAM = 48874;
      end
      6842: begin
        W_PARAM = 16123;
      end
      6843: begin
        W_PARAM = 15831;
      end
      6844: begin
        W_PARAM = 48602;
      end
      6845: begin
        W_PARAM = 15959;
      end
      6846: begin
        W_PARAM = 48969;
      end
      6847: begin
        W_PARAM = 48812;
      end
      6848: begin
        W_PARAM = 16119;
      end
      6849: begin
        W_PARAM = 48814;
      end
      6850: begin
        W_PARAM = 16130;
      end
      6851: begin
        W_PARAM = 48899;
      end
      6852: begin
        W_PARAM = 48790;
      end
      6853: begin
        W_PARAM = 16040;
      end
      6854: begin
        W_PARAM = 48704;
      end
      6855: begin
        W_PARAM = 16161;
      end
      6856: begin
        W_PARAM = 48954;
      end
      6857: begin
        W_PARAM = 16053;
      end
      6858: begin
        W_PARAM = 16062;
      end
      6859: begin
        W_PARAM = 48880;
      end
      6860: begin
        W_PARAM = 16008;
      end
      6861: begin
        W_PARAM = 48814;
      end
      6862: begin
        W_PARAM = 16199;
      end
      6863: begin
        W_PARAM = 16114;
      end
      6864: begin
        W_PARAM = 48761;
      end
      6865: begin
        W_PARAM = 16069;
      end
      6866: begin
        W_PARAM = 48920;
      end
      6867: begin
        W_PARAM = 48731;
      end
      6868: begin
        W_PARAM = 16065;
      end
      6869: begin
        W_PARAM = 48994;
      end
      6870: begin
        W_PARAM = 48622;
      end
      6871: begin
        W_PARAM = 48406;
      end
      6872: begin
        W_PARAM = 48689;
      end
      6873: begin
        W_PARAM = 15981;
      end
      6874: begin
        W_PARAM = 48759;
      end
      6875: begin
        W_PARAM = 16101;
      end
      6876: begin
        W_PARAM = 48777;
      end
      6877: begin
        W_PARAM = 48753;
      end
      6878: begin
        W_PARAM = 15994;
      end
      6879: begin
        W_PARAM = 15896;
      end
      6880: begin
        W_PARAM = 48580;
      end
      6881: begin
        W_PARAM = 49041;
      end
      6882: begin
        W_PARAM = 48676;
      end
      6883: begin
        W_PARAM = 16134;
      end
      6884: begin
        W_PARAM = 15860;
      end
      6885: begin
        W_PARAM = 48403;
      end
      6886: begin
        W_PARAM = 16024;
      end
      6887: begin
        W_PARAM = 48777;
      end
      6888: begin
        W_PARAM = 16253;
      end
      6889: begin
        W_PARAM = 48754;
      end
      6890: begin
        W_PARAM = 15859;
      end
      6891: begin
        W_PARAM = 48467;
      end
      6892: begin
        W_PARAM = 16016;
      end
      6893: begin
        W_PARAM = 16038;
      end
      6894: begin
        W_PARAM = 48792;
      end
      6895: begin
        W_PARAM = 16094;
      end
      6896: begin
        W_PARAM = 15910;
      end
      6897: begin
        W_PARAM = 48583;
      end
      6898: begin
        W_PARAM = 48960;
      end
      6899: begin
        W_PARAM = 48639;
      end
      6900: begin
        W_PARAM = 48770;
      end
      6901: begin
        W_PARAM = 15963;
      end
      6902: begin
        W_PARAM = 16160;
      end
      6903: begin
        W_PARAM = 48920;
      end
      6904: begin
        W_PARAM = 48635;
      end
      6905: begin
        W_PARAM = 16133;
      end
      6906: begin
        W_PARAM = 48595;
      end
      6907: begin
        W_PARAM = 48977;
      end
      6908: begin
        W_PARAM = 16099;
      end
      6909: begin
        W_PARAM = 15784;
      end
      6910: begin
        W_PARAM = 48975;
      end
      6911: begin
        W_PARAM = 16006;
      end
      6912: begin
        W_PARAM = 15754;
      end
      6913: begin
        W_PARAM = 48776;
      end
      6914: begin
        W_PARAM = 15979;
      end
      6915: begin
        W_PARAM = 48563;
      end
      6916: begin
        W_PARAM = 48797;
      end
      6917: begin
        W_PARAM = 48871;
      end
      6918: begin
        W_PARAM = 16293;
      end
      6919: begin
        W_PARAM = 15761;
      end
      6920: begin
        W_PARAM = 48997;
      end
      6921: begin
        W_PARAM = 48471;
      end
      6922: begin
        W_PARAM = 15824;
      end
      6923: begin
        W_PARAM = 15631;
      end
      6924: begin
        W_PARAM = 15889;
      end
      6925: begin
        W_PARAM = 15956;
      end
      6926: begin
        W_PARAM = 48622;
      end
      6927: begin
        W_PARAM = 48661;
      end
      6928: begin
        W_PARAM = 15937;
      end
      6929: begin
        W_PARAM = 16137;
      end
      6930: begin
        W_PARAM = 48931;
      end
      6931: begin
        W_PARAM = 48585;
      end
      6932: begin
        W_PARAM = 16221;
      end
      6933: begin
        W_PARAM = 15916;
      end
      6934: begin
        W_PARAM = 15992;
      end
      6935: begin
        W_PARAM = 48585;
      end
      6936: begin
        W_PARAM = 48667;
      end
      6937: begin
        W_PARAM = 48837;
      end
      6938: begin
        W_PARAM = 48537;
      end
      6939: begin
        W_PARAM = 15920;
      end
      6940: begin
        W_PARAM = 48819;
      end
      6941: begin
        W_PARAM = 48798;
      end
      6942: begin
        W_PARAM = 15664;
      end
      6943: begin
        W_PARAM = 48513;
      end
      6944: begin
        W_PARAM = 15951;
      end
      6945: begin
        W_PARAM = 16152;
      end
      6946: begin
        W_PARAM = 48527;
      end
      6947: begin
        W_PARAM = 48891;
      end
      6948: begin
        W_PARAM = 47737;
      end
      6949: begin
        W_PARAM = 16098;
      end
      6950: begin
        W_PARAM = 48699;
      end
      6951: begin
        W_PARAM = 48603;
      end
      6952: begin
        W_PARAM = 16053;
      end
      6953: begin
        W_PARAM = 48415;
      end
      6954: begin
        W_PARAM = 15432;
      end
      6955: begin
        W_PARAM = 16036;
      end
      6956: begin
        W_PARAM = 48333;
      end
      6957: begin
        W_PARAM = 48972;
      end
      6958: begin
        W_PARAM = 48587;
      end
      6959: begin
        W_PARAM = 16144;
      end
      6960: begin
        W_PARAM = 48271;
      end
      6961: begin
        W_PARAM = 48513;
      end
      6962: begin
        W_PARAM = 16270;
      end
      6963: begin
        W_PARAM = 48619;
      end
      6964: begin
        W_PARAM = 48749;
      end
      6965: begin
        W_PARAM = 15979;
      end
      6966: begin
        W_PARAM = 48006;
      end
      6967: begin
        W_PARAM = 48804;
      end
      6968: begin
        W_PARAM = 48783;
      end
      6969: begin
        W_PARAM = 48798;
      end
      6970: begin
        W_PARAM = 47748;
      end
      6971: begin
        W_PARAM = 15684;
      end
      6972: begin
        W_PARAM = 16156;
      end
      6973: begin
        W_PARAM = 48257;
      end
      6974: begin
        W_PARAM = 15765;
      end
      6975: begin
        W_PARAM = 48697;
      end
      6976: begin
        W_PARAM = 47451;
      end
      6977: begin
        W_PARAM = 48669;
      end
      6978: begin
        W_PARAM = 48641;
      end
      6979: begin
        W_PARAM = 48770;
      end
      6980: begin
        W_PARAM = 46095;
      end
      6981: begin
        W_PARAM = 15397;
      end
      6982: begin
        W_PARAM = 15853;
      end
      6983: begin
        W_PARAM = 46989;
      end
      6984: begin
        W_PARAM = 47422;
      end
      6985: begin
        W_PARAM = 48023;
      end
      6986: begin
        W_PARAM = 47013;
      end
      6987: begin
        W_PARAM = 46466;
      end
      6988: begin
        W_PARAM = 48326;
      end
      6989: begin
        W_PARAM = 48582;
      end
      6990: begin
        W_PARAM = 0;
      end
      6991: begin
        W_PARAM = 0;
      end
      6992: begin
        W_PARAM = 0;
      end
      6993: begin
        W_PARAM = 0;
      end
      6994: begin
        W_PARAM = 0;
      end
      6995: begin
        W_PARAM = 0;
      end
      6996: begin
        W_PARAM = 0;
      end
      6997: begin
        W_PARAM = 0;
      end
      6998: begin
        W_PARAM = 0;
      end
      6999: begin
        W_PARAM = 0;
      end
      7000: begin
        W_PARAM = 0;
      end
      7001: begin
        W_PARAM = 0;
      end
      7002: begin
        W_PARAM = 0;
      end
      7003: begin
        W_PARAM = 0;
      end
      7004: begin
        W_PARAM = 0;
      end
      7005: begin
        W_PARAM = 0;
      end
      7006: begin
        W_PARAM = 0;
      end
      7007: begin
        W_PARAM = 0;
      end
      7008: begin
        W_PARAM = 0;
      end
      7009: begin
        W_PARAM = 0;
      end
      7010: begin
        W_PARAM = 0;
      end
      7011: begin
        W_PARAM = 0;
      end
      7012: begin
        W_PARAM = 0;
      end
      7013: begin
        W_PARAM = 0;
      end
      7014: begin
        W_PARAM = 0;
      end
      7015: begin
        W_PARAM = 0;
      end
      7016: begin
        W_PARAM = 0;
      end
      7017: begin
        W_PARAM = 0;
      end
      7018: begin
        W_PARAM = 0;
      end
      7019: begin
        W_PARAM = 0;
      end
      7020: begin
        W_PARAM = 46989;
      end
      7021: begin
        W_PARAM = 46019;
      end
      7022: begin
        W_PARAM = 47174;
      end
      7023: begin
        W_PARAM = 15401;
      end
      7024: begin
        W_PARAM = 47430;
      end
      7025: begin
        W_PARAM = 46809;
      end
      7026: begin
        W_PARAM = 45973;
      end
      7027: begin
        W_PARAM = 48259;
      end
      7028: begin
        W_PARAM = 47900;
      end
      7029: begin
        W_PARAM = 15369;
      end
      7030: begin
        W_PARAM = 47113;
      end
      7031: begin
        W_PARAM = 48407;
      end
      7032: begin
        W_PARAM = 48484;
      end
      7033: begin
        W_PARAM = 48777;
      end
      7034: begin
        W_PARAM = 46981;
      end
      7035: begin
        W_PARAM = 16010;
      end
      7036: begin
        W_PARAM = 46998;
      end
      7037: begin
        W_PARAM = 15858;
      end
      7038: begin
        W_PARAM = 48082;
      end
      7039: begin
        W_PARAM = 48296;
      end
      7040: begin
        W_PARAM = 47946;
      end
      7041: begin
        W_PARAM = 48682;
      end
      7042: begin
        W_PARAM = 48649;
      end
      7043: begin
        W_PARAM = 48782;
      end
      7044: begin
        W_PARAM = 15678;
      end
      7045: begin
        W_PARAM = 16060;
      end
      7046: begin
        W_PARAM = 47785;
      end
      7047: begin
        W_PARAM = 16053;
      end
      7048: begin
        W_PARAM = 48791;
      end
      7049: begin
        W_PARAM = 15841;
      end
      7050: begin
        W_PARAM = 48529;
      end
      7051: begin
        W_PARAM = 48826;
      end
      7052: begin
        W_PARAM = 48721;
      end
      7053: begin
        W_PARAM = 15915;
      end
      7054: begin
        W_PARAM = 48577;
      end
      7055: begin
        W_PARAM = 15822;
      end
      7056: begin
        W_PARAM = 48027;
      end
      7057: begin
        W_PARAM = 48437;
      end
      7058: begin
        W_PARAM = 48914;
      end
      7059: begin
        W_PARAM = 16267;
      end
      7060: begin
        W_PARAM = 48842;
      end
      7061: begin
        W_PARAM = 48846;
      end
      7062: begin
        W_PARAM = 47882;
      end
      7063: begin
        W_PARAM = 16185;
      end
      7064: begin
        W_PARAM = 48848;
      end
      7065: begin
        W_PARAM = 15824;
      end
      7066: begin
        W_PARAM = 48188;
      end
      7067: begin
        W_PARAM = 48590;
      end
      7068: begin
        W_PARAM = 48640;
      end
      7069: begin
        W_PARAM = 16158;
      end
      7070: begin
        W_PARAM = 48858;
      end
      7071: begin
        W_PARAM = 48900;
      end
      7072: begin
        W_PARAM = 48757;
      end
      7073: begin
        W_PARAM = 16283;
      end
      7074: begin
        W_PARAM = 48877;
      end
      7075: begin
        W_PARAM = 15945;
      end
      7076: begin
        W_PARAM = 48340;
      end
      7077: begin
        W_PARAM = 48288;
      end
      7078: begin
        W_PARAM = 48469;
      end
      7079: begin
        W_PARAM = 16042;
      end
      7080: begin
        W_PARAM = 48899;
      end
      7081: begin
        W_PARAM = 48839;
      end
      7082: begin
        W_PARAM = 48981;
      end
      7083: begin
        W_PARAM = 16356;
      end
      7084: begin
        W_PARAM = 49005;
      end
      7085: begin
        W_PARAM = 15355;
      end
      7086: begin
        W_PARAM = 48585;
      end
      7087: begin
        W_PARAM = 16164;
      end
      7088: begin
        W_PARAM = 48808;
      end
      7089: begin
        W_PARAM = 16167;
      end
      7090: begin
        W_PARAM = 48933;
      end
      7091: begin
        W_PARAM = 48890;
      end
      7092: begin
        W_PARAM = 49048;
      end
      7093: begin
        W_PARAM = 16302;
      end
      7094: begin
        W_PARAM = 48819;
      end
      7095: begin
        W_PARAM = 16145;
      end
      7096: begin
        W_PARAM = 48642;
      end
      7097: begin
        W_PARAM = 16207;
      end
      7098: begin
        W_PARAM = 48825;
      end
      7099: begin
        W_PARAM = 16087;
      end
      7100: begin
        W_PARAM = 49026;
      end
      7101: begin
        W_PARAM = 49088;
      end
      7102: begin
        W_PARAM = 48941;
      end
      7103: begin
        W_PARAM = 16257;
      end
      7104: begin
        W_PARAM = 16004;
      end
      7105: begin
        W_PARAM = 16134;
      end
      7106: begin
        W_PARAM = 48591;
      end
      7107: begin
        W_PARAM = 16008;
      end
      7108: begin
        W_PARAM = 16149;
      end
      7109: begin
        W_PARAM = 16166;
      end
      7110: begin
        W_PARAM = 49002;
      end
      7111: begin
        W_PARAM = 49040;
      end
      7112: begin
        W_PARAM = 48952;
      end
      7113: begin
        W_PARAM = 16137;
      end
      7114: begin
        W_PARAM = 48659;
      end
      7115: begin
        W_PARAM = 16179;
      end
      7116: begin
        W_PARAM = 48482;
      end
      7117: begin
        W_PARAM = 16249;
      end
      7118: begin
        W_PARAM = 16030;
      end
      7119: begin
        W_PARAM = 16098;
      end
      7120: begin
        W_PARAM = 49073;
      end
      7121: begin
        W_PARAM = 48845;
      end
      7122: begin
        W_PARAM = 48731;
      end
      7123: begin
        W_PARAM = 16301;
      end
      7124: begin
        W_PARAM = 48952;
      end
      7125: begin
        W_PARAM = 16148;
      end
      7126: begin
        W_PARAM = 15792;
      end
      7127: begin
        W_PARAM = 16145;
      end
      7128: begin
        W_PARAM = 48792;
      end
      7129: begin
        W_PARAM = 16088;
      end
      7130: begin
        W_PARAM = 49064;
      end
      7131: begin
        W_PARAM = 48862;
      end
      7132: begin
        W_PARAM = 48646;
      end
      7133: begin
        W_PARAM = 16234;
      end
      7134: begin
        W_PARAM = 48568;
      end
      7135: begin
        W_PARAM = 16175;
      end
      7136: begin
        W_PARAM = 48746;
      end
      7137: begin
        W_PARAM = 15988;
      end
      7138: begin
        W_PARAM = 48618;
      end
      7139: begin
        W_PARAM = 16112;
      end
      7140: begin
        W_PARAM = 49069;
      end
      7141: begin
        W_PARAM = 48919;
      end
      7142: begin
        W_PARAM = 15981;
      end
      7143: begin
        W_PARAM = 16143;
      end
      7144: begin
        W_PARAM = 48712;
      end
      7145: begin
        W_PARAM = 48629;
      end
      7146: begin
        W_PARAM = 48771;
      end
      7147: begin
        W_PARAM = 16126;
      end
      7148: begin
        W_PARAM = 16058;
      end
      7149: begin
        W_PARAM = 16222;
      end
      7150: begin
        W_PARAM = 49052;
      end
      7151: begin
        W_PARAM = 48958;
      end
      7152: begin
        W_PARAM = 16138;
      end
      7153: begin
        W_PARAM = 16006;
      end
      7154: begin
        W_PARAM = 48654;
      end
      7155: begin
        W_PARAM = 16227;
      end
      7156: begin
        W_PARAM = 48798;
      end
      7157: begin
        W_PARAM = 16016;
      end
      7158: begin
        W_PARAM = 16079;
      end
      7159: begin
        W_PARAM = 15620;
      end
      7160: begin
        W_PARAM = 48956;
      end
      7161: begin
        W_PARAM = 49040;
      end
      7162: begin
        W_PARAM = 16024;
      end
      7163: begin
        W_PARAM = 16187;
      end
      7164: begin
        W_PARAM = 48881;
      end
      7165: begin
        W_PARAM = 16083;
      end
      7166: begin
        W_PARAM = 48762;
      end
      7167: begin
        W_PARAM = 15932;
      end
      7168: begin
        W_PARAM = 16117;
      end
      7169: begin
        W_PARAM = 16113;
      end
      7170: begin
        W_PARAM = 49039;
      end
      7171: begin
        W_PARAM = 48964;
      end
      7172: begin
        W_PARAM = 15910;
      end
      7173: begin
        W_PARAM = 16157;
      end
      7174: begin
        W_PARAM = 48812;
      end
      7175: begin
        W_PARAM = 16158;
      end
      7176: begin
        W_PARAM = 48649;
      end
      7177: begin
        W_PARAM = 48639;
      end
      7178: begin
        W_PARAM = 16194;
      end
      7179: begin
        W_PARAM = 16039;
      end
      7180: begin
        W_PARAM = 49033;
      end
      7181: begin
        W_PARAM = 48899;
      end
      7182: begin
        W_PARAM = 48915;
      end
      7183: begin
        W_PARAM = 16127;
      end
      7184: begin
        W_PARAM = 48669;
      end
      7185: begin
        W_PARAM = 16143;
      end
      7186: begin
        W_PARAM = 48629;
      end
      7187: begin
        W_PARAM = 16171;
      end
      7188: begin
        W_PARAM = 16034;
      end
      7189: begin
        W_PARAM = 16071;
      end
      7190: begin
        W_PARAM = 48903;
      end
      7191: begin
        W_PARAM = 48885;
      end
      7192: begin
        W_PARAM = 48973;
      end
      7193: begin
        W_PARAM = 16236;
      end
      7194: begin
        W_PARAM = 48971;
      end
      7195: begin
        W_PARAM = 16195;
      end
      7196: begin
        W_PARAM = 48515;
      end
      7197: begin
        W_PARAM = 15963;
      end
      7198: begin
        W_PARAM = 16001;
      end
      7199: begin
        W_PARAM = 16132;
      end
      7200: begin
        W_PARAM = 48924;
      end
      7201: begin
        W_PARAM = 48669;
      end
      7202: begin
        W_PARAM = 48920;
      end
      7203: begin
        W_PARAM = 15880;
      end
      7204: begin
        W_PARAM = 48858;
      end
      7205: begin
        W_PARAM = 16154;
      end
      7206: begin
        W_PARAM = 48410;
      end
      7207: begin
        W_PARAM = 48444;
      end
      7208: begin
        W_PARAM = 15929;
      end
      7209: begin
        W_PARAM = 16243;
      end
      7210: begin
        W_PARAM = 48868;
      end
      7211: begin
        W_PARAM = 48318;
      end
      7212: begin
        W_PARAM = 48906;
      end
      7213: begin
        W_PARAM = 48871;
      end
      7214: begin
        W_PARAM = 48898;
      end
      7215: begin
        W_PARAM = 16227;
      end
      7216: begin
        W_PARAM = 48287;
      end
      7217: begin
        W_PARAM = 15858;
      end
      7218: begin
        W_PARAM = 48352;
      end
      7219: begin
        W_PARAM = 16257;
      end
      7220: begin
        W_PARAM = 48758;
      end
      7221: begin
        W_PARAM = 48203;
      end
      7222: begin
        W_PARAM = 48906;
      end
      7223: begin
        W_PARAM = 48680;
      end
      7224: begin
        W_PARAM = 48775;
      end
      7225: begin
        W_PARAM = 16261;
      end
      7226: begin
        W_PARAM = 48151;
      end
      7227: begin
        W_PARAM = 16029;
      end
      7228: begin
        W_PARAM = 48617;
      end
      7229: begin
        W_PARAM = 47946;
      end
      7230: begin
        W_PARAM = 48541;
      end
      7231: begin
        W_PARAM = 47683;
      end
      7232: begin
        W_PARAM = 48768;
      end
      7233: begin
        W_PARAM = 48257;
      end
      7234: begin
        W_PARAM = 48781;
      end
      7235: begin
        W_PARAM = 16182;
      end
      7236: begin
        W_PARAM = 47990;
      end
      7237: begin
        W_PARAM = 48625;
      end
      7238: begin
        W_PARAM = 48445;
      end
      7239: begin
        W_PARAM = 15771;
      end
      7240: begin
        W_PARAM = 48119;
      end
      7241: begin
        W_PARAM = 46732;
      end
      7242: begin
        W_PARAM = 48148;
      end
      7243: begin
        W_PARAM = 47372;
      end
      7244: begin
        W_PARAM = 48700;
      end
      7245: begin
        W_PARAM = 16096;
      end
      7246: begin
        W_PARAM = 47544;
      end
      7247: begin
        W_PARAM = 48117;
      end
      7248: begin
        W_PARAM = 48160;
      end
      7249: begin
        W_PARAM = 48737;
      end
      7250: begin
        W_PARAM = 46106;
      end
      7251: begin
        W_PARAM = 46924;
      end
      7252: begin
        W_PARAM = 15826;
      end
      7253: begin
        W_PARAM = 47747;
      end
      7254: begin
        W_PARAM = 47767;
      end
      7255: begin
        W_PARAM = 46863;
      end
      7256: begin
        W_PARAM = 46927;
      end
      7257: begin
        W_PARAM = 48045;
      end
      7258: begin
        W_PARAM = 48278;
      end
      7259: begin
        W_PARAM = 48541;
      end
      7260: begin
        W_PARAM = 46100;
      end
      7261: begin
        W_PARAM = 46964;
      end
      7262: begin
        W_PARAM = 15867;
      end
      7263: begin
        W_PARAM = 46336;
      end
      7264: begin
        W_PARAM = 47434;
      end
      7265: begin
        W_PARAM = 46780;
      end
      7266: begin
        W_PARAM = 46967;
      end
      7267: begin
        W_PARAM = 46457;
      end
      7268: begin
        W_PARAM = 48290;
      end
      7269: begin
        W_PARAM = 48594;
      end
      7270: begin
        W_PARAM = 0;
      end
      7271: begin
        W_PARAM = 0;
      end
      7272: begin
        W_PARAM = 0;
      end
      7273: begin
        W_PARAM = 0;
      end
      7274: begin
        W_PARAM = 0;
      end
      7275: begin
        W_PARAM = 0;
      end
      7276: begin
        W_PARAM = 0;
      end
      7277: begin
        W_PARAM = 0;
      end
      7278: begin
        W_PARAM = 0;
      end
      7279: begin
        W_PARAM = 0;
      end
      7280: begin
        W_PARAM = 0;
      end
      7281: begin
        W_PARAM = 0;
      end
      7282: begin
        W_PARAM = 0;
      end
      7283: begin
        W_PARAM = 0;
      end
      7284: begin
        W_PARAM = 0;
      end
      7285: begin
        W_PARAM = 0;
      end
      7286: begin
        W_PARAM = 0;
      end
      7287: begin
        W_PARAM = 0;
      end
      7288: begin
        W_PARAM = 0;
      end
      7289: begin
        W_PARAM = 0;
      end
      7290: begin
        W_PARAM = 0;
      end
      7291: begin
        W_PARAM = 0;
      end
      7292: begin
        W_PARAM = 0;
      end
      7293: begin
        W_PARAM = 0;
      end
      7294: begin
        W_PARAM = 0;
      end
      7295: begin
        W_PARAM = 0;
      end
      7296: begin
        W_PARAM = 0;
      end
      7297: begin
        W_PARAM = 0;
      end
      7298: begin
        W_PARAM = 0;
      end
      7299: begin
        W_PARAM = 0;
      end
      7300: begin
        W_PARAM = 0;
      end
      7301: begin
        W_PARAM = 0;
      end
      7302: begin
        W_PARAM = 0;
      end
      7303: begin
        W_PARAM = 0;
      end
      7304: begin
        W_PARAM = 0;
      end
      7305: begin
        W_PARAM = 0;
      end
      7306: begin
        W_PARAM = 0;
      end
      7307: begin
        W_PARAM = 0;
      end
      7308: begin
        W_PARAM = 0;
      end
      7309: begin
        W_PARAM = 0;
      end
      7310: begin
        W_PARAM = 0;
      end
      7311: begin
        W_PARAM = 0;
      end
      7312: begin
        W_PARAM = 0;
      end
      7313: begin
        W_PARAM = 0;
      end
      7314: begin
        W_PARAM = 0;
      end
      7315: begin
        W_PARAM = 0;
      end
      7316: begin
        W_PARAM = 0;
      end
      7317: begin
        W_PARAM = 0;
      end
      7318: begin
        W_PARAM = 0;
      end
      7319: begin
        W_PARAM = 0;
      end
      7320: begin
        W_PARAM = 47795;
      end
      7321: begin
        W_PARAM = 47712;
      end
      7322: begin
        W_PARAM = 47638;
      end
      7323: begin
        W_PARAM = 15253;
      end
      7324: begin
        W_PARAM = 15657;
      end
      7325: begin
        W_PARAM = 47919;
      end
      7326: begin
        W_PARAM = 47647;
      end
      7327: begin
        W_PARAM = 48796;
      end
      7328: begin
        W_PARAM = 48281;
      end
      7329: begin
        W_PARAM = 16017;
      end
      7330: begin
        W_PARAM = 48147;
      end
      7331: begin
        W_PARAM = 47948;
      end
      7332: begin
        W_PARAM = 47993;
      end
      7333: begin
        W_PARAM = 15857;
      end
      7334: begin
        W_PARAM = 15772;
      end
      7335: begin
        W_PARAM = 48154;
      end
      7336: begin
        W_PARAM = 47897;
      end
      7337: begin
        W_PARAM = 48929;
      end
      7338: begin
        W_PARAM = 48626;
      end
      7339: begin
        W_PARAM = 16149;
      end
      7340: begin
        W_PARAM = 48513;
      end
      7341: begin
        W_PARAM = 48236;
      end
      7342: begin
        W_PARAM = 48327;
      end
      7343: begin
        W_PARAM = 15943;
      end
      7344: begin
        W_PARAM = 48648;
      end
      7345: begin
        W_PARAM = 48714;
      end
      7346: begin
        W_PARAM = 48111;
      end
      7347: begin
        W_PARAM = 48812;
      end
      7348: begin
        W_PARAM = 48770;
      end
      7349: begin
        W_PARAM = 16213;
      end
      7350: begin
        W_PARAM = 48621;
      end
      7351: begin
        W_PARAM = 48337;
      end
      7352: begin
        W_PARAM = 48532;
      end
      7353: begin
        W_PARAM = 15968;
      end
      7354: begin
        W_PARAM = 48875;
      end
      7355: begin
        W_PARAM = 48919;
      end
      7356: begin
        W_PARAM = 48142;
      end
      7357: begin
        W_PARAM = 15994;
      end
      7358: begin
        W_PARAM = 48396;
      end
      7359: begin
        W_PARAM = 16216;
      end
      7360: begin
        W_PARAM = 48642;
      end
      7361: begin
        W_PARAM = 48407;
      end
      7362: begin
        W_PARAM = 48557;
      end
      7363: begin
        W_PARAM = 15816;
      end
      7364: begin
        W_PARAM = 48918;
      end
      7365: begin
        W_PARAM = 48958;
      end
      7366: begin
        W_PARAM = 48246;
      end
      7367: begin
        W_PARAM = 16070;
      end
      7368: begin
        W_PARAM = 15774;
      end
      7369: begin
        W_PARAM = 16260;
      end
      7370: begin
        W_PARAM = 48770;
      end
      7371: begin
        W_PARAM = 48494;
      end
      7372: begin
        W_PARAM = 48626;
      end
      7373: begin
        W_PARAM = 15633;
      end
      7374: begin
        W_PARAM = 49013;
      end
      7375: begin
        W_PARAM = 48885;
      end
      7376: begin
        W_PARAM = 48408;
      end
      7377: begin
        W_PARAM = 16203;
      end
      7378: begin
        W_PARAM = 48662;
      end
      7379: begin
        W_PARAM = 16284;
      end
      7380: begin
        W_PARAM = 48734;
      end
      7381: begin
        W_PARAM = 48783;
      end
      7382: begin
        W_PARAM = 48519;
      end
      7383: begin
        W_PARAM = 16031;
      end
      7384: begin
        W_PARAM = 49002;
      end
      7385: begin
        W_PARAM = 48606;
      end
      7386: begin
        W_PARAM = 48392;
      end
      7387: begin
        W_PARAM = 16172;
      end
      7388: begin
        W_PARAM = 48869;
      end
      7389: begin
        W_PARAM = 16267;
      end
      7390: begin
        W_PARAM = 48635;
      end
      7391: begin
        W_PARAM = 48765;
      end
      7392: begin
        W_PARAM = 48786;
      end
      7393: begin
        W_PARAM = 16084;
      end
      7394: begin
        W_PARAM = 49043;
      end
      7395: begin
        W_PARAM = 16123;
      end
      7396: begin
        W_PARAM = 48259;
      end
      7397: begin
        W_PARAM = 16058;
      end
      7398: begin
        W_PARAM = 48673;
      end
      7399: begin
        W_PARAM = 16181;
      end
      7400: begin
        W_PARAM = 48487;
      end
      7401: begin
        W_PARAM = 48847;
      end
      7402: begin
        W_PARAM = 48629;
      end
      7403: begin
        W_PARAM = 15943;
      end
      7404: begin
        W_PARAM = 49031;
      end
      7405: begin
        W_PARAM = 16095;
      end
      7406: begin
        W_PARAM = 48225;
      end
      7407: begin
        W_PARAM = 15571;
      end
      7408: begin
        W_PARAM = 48550;
      end
      7409: begin
        W_PARAM = 16265;
      end
      7410: begin
        W_PARAM = 48711;
      end
      7411: begin
        W_PARAM = 48916;
      end
      7412: begin
        W_PARAM = 48787;
      end
      7413: begin
        W_PARAM = 16020;
      end
      7414: begin
        W_PARAM = 49048;
      end
      7415: begin
        W_PARAM = 15999;
      end
      7416: begin
        W_PARAM = 48474;
      end
      7417: begin
        W_PARAM = 16213;
      end
      7418: begin
        W_PARAM = 48436;
      end
      7419: begin
        W_PARAM = 16248;
      end
      7420: begin
        W_PARAM = 48789;
      end
      7421: begin
        W_PARAM = 48830;
      end
      7422: begin
        W_PARAM = 48720;
      end
      7423: begin
        W_PARAM = 16022;
      end
      7424: begin
        W_PARAM = 49098;
      end
      7425: begin
        W_PARAM = 15975;
      end
      7426: begin
        W_PARAM = 48461;
      end
      7427: begin
        W_PARAM = 16208;
      end
      7428: begin
        W_PARAM = 48837;
      end
      7429: begin
        W_PARAM = 16326;
      end
      7430: begin
        W_PARAM = 48737;
      end
      7431: begin
        W_PARAM = 48616;
      end
      7432: begin
        W_PARAM = 48767;
      end
      7433: begin
        W_PARAM = 16024;
      end
      7434: begin
        W_PARAM = 49073;
      end
      7435: begin
        W_PARAM = 16178;
      end
      7436: begin
        W_PARAM = 48376;
      end
      7437: begin
        W_PARAM = 16257;
      end
      7438: begin
        W_PARAM = 48968;
      end
      7439: begin
        W_PARAM = 16198;
      end
      7440: begin
        W_PARAM = 48671;
      end
      7441: begin
        W_PARAM = 48662;
      end
      7442: begin
        W_PARAM = 48812;
      end
      7443: begin
        W_PARAM = 16171;
      end
      7444: begin
        W_PARAM = 49053;
      end
      7445: begin
        W_PARAM = 15964;
      end
      7446: begin
        W_PARAM = 48290;
      end
      7447: begin
        W_PARAM = 16146;
      end
      7448: begin
        W_PARAM = 48890;
      end
      7449: begin
        W_PARAM = 16235;
      end
      7450: begin
        W_PARAM = 48805;
      end
      7451: begin
        W_PARAM = 48632;
      end
      7452: begin
        W_PARAM = 48847;
      end
      7453: begin
        W_PARAM = 16154;
      end
      7454: begin
        W_PARAM = 49050;
      end
      7455: begin
        W_PARAM = 48595;
      end
      7456: begin
        W_PARAM = 48320;
      end
      7457: begin
        W_PARAM = 16214;
      end
      7458: begin
        W_PARAM = 48647;
      end
      7459: begin
        W_PARAM = 16223;
      end
      7460: begin
        W_PARAM = 48725;
      end
      7461: begin
        W_PARAM = 48767;
      end
      7462: begin
        W_PARAM = 48738;
      end
      7463: begin
        W_PARAM = 16051;
      end
      7464: begin
        W_PARAM = 49065;
      end
      7465: begin
        W_PARAM = 48739;
      end
      7466: begin
        W_PARAM = 48316;
      end
      7467: begin
        W_PARAM = 16191;
      end
      7468: begin
        W_PARAM = 48591;
      end
      7469: begin
        W_PARAM = 16288;
      end
      7470: begin
        W_PARAM = 48272;
      end
      7471: begin
        W_PARAM = 48658;
      end
      7472: begin
        W_PARAM = 48439;
      end
      7473: begin
        W_PARAM = 15914;
      end
      7474: begin
        W_PARAM = 49037;
      end
      7475: begin
        W_PARAM = 15781;
      end
      7476: begin
        W_PARAM = 48178;
      end
      7477: begin
        W_PARAM = 16188;
      end
      7478: begin
        W_PARAM = 48807;
      end
      7479: begin
        W_PARAM = 16168;
      end
      7480: begin
        W_PARAM = 48710;
      end
      7481: begin
        W_PARAM = 48388;
      end
      7482: begin
        W_PARAM = 48511;
      end
      7483: begin
        W_PARAM = 15410;
      end
      7484: begin
        W_PARAM = 48928;
      end
      7485: begin
        W_PARAM = 16003;
      end
      7486: begin
        W_PARAM = 47963;
      end
      7487: begin
        W_PARAM = 15659;
      end
      7488: begin
        W_PARAM = 48660;
      end
      7489: begin
        W_PARAM = 16193;
      end
      7490: begin
        W_PARAM = 48751;
      end
      7491: begin
        W_PARAM = 48277;
      end
      7492: begin
        W_PARAM = 48572;
      end
      7493: begin
        W_PARAM = 48291;
      end
      7494: begin
        W_PARAM = 48838;
      end
      7495: begin
        W_PARAM = 15954;
      end
      7496: begin
        W_PARAM = 47928;
      end
      7497: begin
        W_PARAM = 48268;
      end
      7498: begin
        W_PARAM = 48321;
      end
      7499: begin
        W_PARAM = 16151;
      end
      7500: begin
        W_PARAM = 48663;
      end
      7501: begin
        W_PARAM = 47932;
      end
      7502: begin
        W_PARAM = 48408;
      end
      7503: begin
        W_PARAM = 15279;
      end
      7504: begin
        W_PARAM = 48797;
      end
      7505: begin
        W_PARAM = 15788;
      end
      7506: begin
        W_PARAM = 47505;
      end
      7507: begin
        W_PARAM = 16031;
      end
      7508: begin
        W_PARAM = 48002;
      end
      7509: begin
        W_PARAM = 15818;
      end
      7510: begin
        W_PARAM = 48072;
      end
      7511: begin
        W_PARAM = 46648;
      end
      7512: begin
        W_PARAM = 47343;
      end
      7513: begin
        W_PARAM = 47869;
      end
      7514: begin
        W_PARAM = 48442;
      end
      7515: begin
        W_PARAM = 15008;
      end
      7516: begin
        W_PARAM = 46983;
      end
      7517: begin
        W_PARAM = 15446;
      end
      7518: begin
        W_PARAM = 47560;
      end
      7519: begin
        W_PARAM = 15650;
      end
      7520: begin
        W_PARAM = 46851;
      end
      7521: begin
        W_PARAM = 44930;
      end
      7522: begin
        W_PARAM = 46389;
      end
      7523: begin
        W_PARAM = 46062;
      end
      7524: begin
        W_PARAM = 48131;
      end
      7525: begin
        W_PARAM = 47551;
      end
      7526: begin
        W_PARAM = 46440;
      end
      7527: begin
        W_PARAM = 47643;
      end
      7528: begin
        W_PARAM = 46930;
      end
      7529: begin
        W_PARAM = 15379;
      end
      7530: begin
        W_PARAM = 45993;
      end
      7531: begin
        W_PARAM = 45337;
      end
      7532: begin
        W_PARAM = 46383;
      end
      7533: begin
        W_PARAM = 46139;
      end
      7534: begin
        W_PARAM = 45552;
      end
      7535: begin
        W_PARAM = 45540;
      end
      7536: begin
        W_PARAM = 43785;
      end
      7537: begin
        W_PARAM = 14391;
      end
      7538: begin
        W_PARAM = 45979;
      end
      7539: begin
        W_PARAM = 47154;
      end
      7540: begin
        W_PARAM = 0;
      end
      7541: begin
        W_PARAM = 0;
      end
      7542: begin
        W_PARAM = 0;
      end
      7543: begin
        W_PARAM = 0;
      end
      7544: begin
        W_PARAM = 0;
      end
      7545: begin
        W_PARAM = 0;
      end
      7546: begin
        W_PARAM = 0;
      end
      7547: begin
        W_PARAM = 0;
      end
      7548: begin
        W_PARAM = 0;
      end
      7549: begin
        W_PARAM = 0;
      end
      7550: begin
        W_PARAM = 0;
      end
      7551: begin
        W_PARAM = 0;
      end
      7552: begin
        W_PARAM = 0;
      end
      7553: begin
        W_PARAM = 0;
      end
      7554: begin
        W_PARAM = 0;
      end
      7555: begin
        W_PARAM = 0;
      end
      7556: begin
        W_PARAM = 0;
      end
      7557: begin
        W_PARAM = 0;
      end
      7558: begin
        W_PARAM = 0;
      end
      7559: begin
        W_PARAM = 0;
      end
      7560: begin
        W_PARAM = 0;
      end
      7561: begin
        W_PARAM = 0;
      end
      7562: begin
        W_PARAM = 0;
      end
      7563: begin
        W_PARAM = 0;
      end
      7564: begin
        W_PARAM = 0;
      end
      7565: begin
        W_PARAM = 0;
      end
      7566: begin
        W_PARAM = 0;
      end
      7567: begin
        W_PARAM = 0;
      end
      7568: begin
        W_PARAM = 0;
      end
      7569: begin
        W_PARAM = 0;
      end
      7570: begin
        W_PARAM = 0;
      end
      7571: begin
        W_PARAM = 0;
      end
      7572: begin
        W_PARAM = 0;
      end
      7573: begin
        W_PARAM = 0;
      end
      7574: begin
        W_PARAM = 0;
      end
      7575: begin
        W_PARAM = 0;
      end
      7576: begin
        W_PARAM = 0;
      end
      7577: begin
        W_PARAM = 0;
      end
      7578: begin
        W_PARAM = 0;
      end
      7579: begin
        W_PARAM = 0;
      end
      7580: begin
        W_PARAM = 0;
      end
      7581: begin
        W_PARAM = 0;
      end
      7582: begin
        W_PARAM = 0;
      end
      7583: begin
        W_PARAM = 0;
      end
      7584: begin
        W_PARAM = 0;
      end
      7585: begin
        W_PARAM = 0;
      end
      7586: begin
        W_PARAM = 0;
      end
      7587: begin
        W_PARAM = 0;
      end
      7588: begin
        W_PARAM = 0;
      end
      7589: begin
        W_PARAM = 0;
      end
      7590: begin
        W_PARAM = 0;
      end
      7591: begin
        W_PARAM = 0;
      end
      7592: begin
        W_PARAM = 0;
      end
      7593: begin
        W_PARAM = 0;
      end
      7594: begin
        W_PARAM = 0;
      end
      7595: begin
        W_PARAM = 0;
      end
      7596: begin
        W_PARAM = 0;
      end
      7597: begin
        W_PARAM = 0;
      end
      7598: begin
        W_PARAM = 0;
      end
      7599: begin
        W_PARAM = 0;
      end
      7600: begin
        W_PARAM = 46350;
      end
      7601: begin
        W_PARAM = 46389;
      end
      7602: begin
        W_PARAM = 45961;
      end
      7603: begin
        W_PARAM = 46359;
      end
      7604: begin
        W_PARAM = 45718;
      end
      7605: begin
        W_PARAM = 45985;
      end
      7606: begin
        W_PARAM = 44463;
      end
      7607: begin
        W_PARAM = 15077;
      end
      7608: begin
        W_PARAM = 46856;
      end
      7609: begin
        W_PARAM = 47844;
      end
      7610: begin
        W_PARAM = 46898;
      end
      7611: begin
        W_PARAM = 46563;
      end
      7612: begin
        W_PARAM = 46601;
      end
      7613: begin
        W_PARAM = 46545;
      end
      7614: begin
        W_PARAM = 46131;
      end
      7615: begin
        W_PARAM = 46538;
      end
      7616: begin
        W_PARAM = 45008;
      end
      7617: begin
        W_PARAM = 15278;
      end
      7618: begin
        W_PARAM = 47033;
      end
      7619: begin
        W_PARAM = 48044;
      end
      7620: begin
        W_PARAM = 47106;
      end
      7621: begin
        W_PARAM = 46537;
      end
      7622: begin
        W_PARAM = 46894;
      end
      7623: begin
        W_PARAM = 47167;
      end
      7624: begin
        W_PARAM = 48399;
      end
      7625: begin
        W_PARAM = 47253;
      end
      7626: begin
        W_PARAM = 46181;
      end
      7627: begin
        W_PARAM = 47986;
      end
      7628: begin
        W_PARAM = 47225;
      end
      7629: begin
        W_PARAM = 15647;
      end
      7630: begin
        W_PARAM = 47402;
      end
      7631: begin
        W_PARAM = 46575;
      end
      7632: begin
        W_PARAM = 47210;
      end
      7633: begin
        W_PARAM = 47329;
      end
      7634: begin
        W_PARAM = 48715;
      end
      7635: begin
        W_PARAM = 47639;
      end
      7636: begin
        W_PARAM = 47714;
      end
      7637: begin
        W_PARAM = 48387;
      end
      7638: begin
        W_PARAM = 47481;
      end
      7639: begin
        W_PARAM = 15981;
      end
      7640: begin
        W_PARAM = 47801;
      end
      7641: begin
        W_PARAM = 47567;
      end
      7642: begin
        W_PARAM = 47610;
      end
      7643: begin
        W_PARAM = 47644;
      end
      7644: begin
        W_PARAM = 48708;
      end
      7645: begin
        W_PARAM = 47795;
      end
      7646: begin
        W_PARAM = 48015;
      end
      7647: begin
        W_PARAM = 15510;
      end
      7648: begin
        W_PARAM = 47715;
      end
      7649: begin
        W_PARAM = 15931;
      end
      7650: begin
        W_PARAM = 47915;
      end
      7651: begin
        W_PARAM = 47704;
      end
      7652: begin
        W_PARAM = 47750;
      end
      7653: begin
        W_PARAM = 47957;
      end
      7654: begin
        W_PARAM = 48506;
      end
      7655: begin
        W_PARAM = 47794;
      end
      7656: begin
        W_PARAM = 47998;
      end
      7657: begin
        W_PARAM = 15361;
      end
      7658: begin
        W_PARAM = 47880;
      end
      7659: begin
        W_PARAM = 15755;
      end
      7660: begin
        W_PARAM = 47875;
      end
      7661: begin
        W_PARAM = 48087;
      end
      7662: begin
        W_PARAM = 48278;
      end
      7663: begin
        W_PARAM = 48319;
      end
      7664: begin
        W_PARAM = 48702;
      end
      7665: begin
        W_PARAM = 15490;
      end
      7666: begin
        W_PARAM = 47802;
      end
      7667: begin
        W_PARAM = 15981;
      end
      7668: begin
        W_PARAM = 48480;
      end
      7669: begin
        W_PARAM = 15670;
      end
      7670: begin
        W_PARAM = 47955;
      end
      7671: begin
        W_PARAM = 48021;
      end
      7672: begin
        W_PARAM = 48138;
      end
      7673: begin
        W_PARAM = 48226;
      end
      7674: begin
        W_PARAM = 48617;
      end
      7675: begin
        W_PARAM = 15642;
      end
      7676: begin
        W_PARAM = 47872;
      end
      7677: begin
        W_PARAM = 15753;
      end
      7678: begin
        W_PARAM = 48165;
      end
      7679: begin
        W_PARAM = 15699;
      end
      7680: begin
        W_PARAM = 47907;
      end
      7681: begin
        W_PARAM = 48204;
      end
      7682: begin
        W_PARAM = 47853;
      end
      7683: begin
        W_PARAM = 48184;
      end
      7684: begin
        W_PARAM = 48637;
      end
      7685: begin
        W_PARAM = 15617;
      end
      7686: begin
        W_PARAM = 47812;
      end
      7687: begin
        W_PARAM = 15619;
      end
      7688: begin
        W_PARAM = 48435;
      end
      7689: begin
        W_PARAM = 15880;
      end
      7690: begin
        W_PARAM = 48030;
      end
      7691: begin
        W_PARAM = 48192;
      end
      7692: begin
        W_PARAM = 47893;
      end
      7693: begin
        W_PARAM = 48207;
      end
      7694: begin
        W_PARAM = 48556;
      end
      7695: begin
        W_PARAM = 15218;
      end
      7696: begin
        W_PARAM = 47963;
      end
      7697: begin
        W_PARAM = 16134;
      end
      7698: begin
        W_PARAM = 48399;
      end
      7699: begin
        W_PARAM = 48831;
      end
      7700: begin
        W_PARAM = 48147;
      end
      7701: begin
        W_PARAM = 48051;
      end
      7702: begin
        W_PARAM = 47819;
      end
      7703: begin
        W_PARAM = 48214;
      end
      7704: begin
        W_PARAM = 48847;
      end
      7705: begin
        W_PARAM = 48298;
      end
      7706: begin
        W_PARAM = 47904;
      end
      7707: begin
        W_PARAM = 16059;
      end
      7708: begin
        W_PARAM = 48139;
      end
      7709: begin
        W_PARAM = 15820;
      end
      7710: begin
        W_PARAM = 48250;
      end
      7711: begin
        W_PARAM = 47752;
      end
      7712: begin
        W_PARAM = 47798;
      end
      7713: begin
        W_PARAM = 48139;
      end
      7714: begin
        W_PARAM = 48728;
      end
      7715: begin
        W_PARAM = 48257;
      end
      7716: begin
        W_PARAM = 47730;
      end
      7717: begin
        W_PARAM = 16051;
      end
      7718: begin
        W_PARAM = 48158;
      end
      7719: begin
        W_PARAM = 48563;
      end
      7720: begin
        W_PARAM = 48168;
      end
      7721: begin
        W_PARAM = 47747;
      end
      7722: begin
        W_PARAM = 47802;
      end
      7723: begin
        W_PARAM = 48294;
      end
      7724: begin
        W_PARAM = 48561;
      end
      7725: begin
        W_PARAM = 48252;
      end
      7726: begin
        W_PARAM = 47739;
      end
      7727: begin
        W_PARAM = 15961;
      end
      7728: begin
        W_PARAM = 48068;
      end
      7729: begin
        W_PARAM = 48528;
      end
      7730: begin
        W_PARAM = 47846;
      end
      7731: begin
        W_PARAM = 48415;
      end
      7732: begin
        W_PARAM = 47774;
      end
      7733: begin
        W_PARAM = 48199;
      end
      7734: begin
        W_PARAM = 48503;
      end
      7735: begin
        W_PARAM = 48212;
      end
      7736: begin
        W_PARAM = 47438;
      end
      7737: begin
        W_PARAM = 16047;
      end
      7738: begin
        W_PARAM = 48054;
      end
      7739: begin
        W_PARAM = 48726;
      end
      7740: begin
        W_PARAM = 48091;
      end
      7741: begin
        W_PARAM = 48640;
      end
      7742: begin
        W_PARAM = 47629;
      end
      7743: begin
        W_PARAM = 48043;
      end
      7744: begin
        W_PARAM = 48541;
      end
      7745: begin
        W_PARAM = 48148;
      end
      7746: begin
        W_PARAM = 47079;
      end
      7747: begin
        W_PARAM = 16054;
      end
      7748: begin
        W_PARAM = 48019;
      end
      7749: begin
        W_PARAM = 48644;
      end
      7750: begin
        W_PARAM = 48085;
      end
      7751: begin
        W_PARAM = 47792;
      end
      7752: begin
        W_PARAM = 47486;
      end
      7753: begin
        W_PARAM = 48045;
      end
      7754: begin
        W_PARAM = 48545;
      end
      7755: begin
        W_PARAM = 48296;
      end
      7756: begin
        W_PARAM = 46742;
      end
      7757: begin
        W_PARAM = 16050;
      end
      7758: begin
        W_PARAM = 47940;
      end
      7759: begin
        W_PARAM = 48750;
      end
      7760: begin
        W_PARAM = 47921;
      end
      7761: begin
        W_PARAM = 47040;
      end
      7762: begin
        W_PARAM = 48166;
      end
      7763: begin
        W_PARAM = 47915;
      end
      7764: begin
        W_PARAM = 48117;
      end
      7765: begin
        W_PARAM = 48549;
      end
      7766: begin
        W_PARAM = 46848;
      end
      7767: begin
        W_PARAM = 15869;
      end
      7768: begin
        W_PARAM = 47989;
      end
      7769: begin
        W_PARAM = 48262;
      end
      7770: begin
        W_PARAM = 48471;
      end
      7771: begin
        W_PARAM = 46765;
      end
      7772: begin
        W_PARAM = 48142;
      end
      7773: begin
        W_PARAM = 47542;
      end
      7774: begin
        W_PARAM = 48347;
      end
      7775: begin
        W_PARAM = 48423;
      end
      7776: begin
        W_PARAM = 46973;
      end
      7777: begin
        W_PARAM = 15764;
      end
      7778: begin
        W_PARAM = 47846;
      end
      7779: begin
        W_PARAM = 15727;
      end
      7780: begin
        W_PARAM = 48683;
      end
      7781: begin
        W_PARAM = 46726;
      end
      7782: begin
        W_PARAM = 48411;
      end
      7783: begin
        W_PARAM = 47496;
      end
      7784: begin
        W_PARAM = 48561;
      end
      7785: begin
        W_PARAM = 48306;
      end
      7786: begin
        W_PARAM = 47156;
      end
      7787: begin
        W_PARAM = 15986;
      end
      7788: begin
        W_PARAM = 47820;
      end
      7789: begin
        W_PARAM = 15777;
      end
      7790: begin
        W_PARAM = 48412;
      end
      7791: begin
        W_PARAM = 46448;
      end
      7792: begin
        W_PARAM = 47650;
      end
      7793: begin
        W_PARAM = 46780;
      end
      7794: begin
        W_PARAM = 48292;
      end
      7795: begin
        W_PARAM = 48035;
      end
      7796: begin
        W_PARAM = 46885;
      end
      7797: begin
        W_PARAM = 15813;
      end
      7798: begin
        W_PARAM = 47539;
      end
      7799: begin
        W_PARAM = 48387;
      end
      7800: begin
        W_PARAM = 0;
      end
      7801: begin
        W_PARAM = 0;
      end
      7802: begin
        W_PARAM = 0;
      end
      7803: begin
        W_PARAM = 0;
      end
      7804: begin
        W_PARAM = 0;
      end
      7805: begin
        W_PARAM = 0;
      end
      7806: begin
        W_PARAM = 0;
      end
      7807: begin
        W_PARAM = 0;
      end
      7808: begin
        W_PARAM = 0;
      end
      7809: begin
        W_PARAM = 0;
      end
      7810: begin
        W_PARAM = 0;
      end
      7811: begin
        W_PARAM = 0;
      end
      7812: begin
        W_PARAM = 0;
      end
      7813: begin
        W_PARAM = 0;
      end
      7814: begin
        W_PARAM = 0;
      end
      7815: begin
        W_PARAM = 0;
      end
      7816: begin
        W_PARAM = 0;
      end
      7817: begin
        W_PARAM = 0;
      end
      7818: begin
        W_PARAM = 0;
      end
      7819: begin
        W_PARAM = 0;
      end
      7820: begin
        W_PARAM = 0;
      end
      7821: begin
        W_PARAM = 0;
      end
      7822: begin
        W_PARAM = 0;
      end
      7823: begin
        W_PARAM = 0;
      end
      7824: begin
        W_PARAM = 0;
      end
      7825: begin
        W_PARAM = 0;
      end
      7826: begin
        W_PARAM = 0;
      end
      7827: begin
        W_PARAM = 0;
      end
      7828: begin
        W_PARAM = 0;
      end
      7829: begin
        W_PARAM = 0;
      end
      7830: begin
        W_PARAM = 0;
      end
      7831: begin
        W_PARAM = 0;
      end
      7832: begin
        W_PARAM = 0;
      end
      7833: begin
        W_PARAM = 0;
      end
      7834: begin
        W_PARAM = 0;
      end
      7835: begin
        W_PARAM = 0;
      end
      7836: begin
        W_PARAM = 0;
      end
      7837: begin
        W_PARAM = 0;
      end
      7838: begin
        W_PARAM = 0;
      end
      7839: begin
        W_PARAM = 0;
      end
    endcase
  end
  endfunction
  assign i3 = (i2 + 1);
  assign i_inl1_inl24 = (i_inl1_inl23 + 1);
  assign i_inl1_inl2_inl15 = (i_inl1_inl2_inl14 + 1);
  assign i_inl2_inl24 = (i_inl2_inl23 + 1);
  assign i_inl2_inl2_inl15 = (i_inl2_inl2_inl14 + 1);
  assign j4 = (j3 + 1);
  assign j7 = (j6 + 1);
  assign mul_result1_inl16 = c1196 ? 0 : (c1197 && c1200) ? 0 : (c1197 && (c1205 || c1204)) ? x_w_inl1_inl1 : 'bz;
  assign new_b_n_inl2 = (t572_inl2 + t575_inl2);
  assign new_b_n_inl2_inl1 = (t572_inl2_inl1 + t575_inl2_inl1);
  assign new_n_inl1_inl14 = (new_n_inl1_inl13 >>> 8);
  assign new_n_inl1_inl15 = (new_n_inl1_inl13 >>> 7);
  assign new_n_inl1_inl16 = c1204 ? new_n_inl1_inl14 : c1205 ? new_n_inl1_inl15 : 'bz;
  assign new_n_inl1_inl17 = (new_n_inl1_inl16 & 127);
  assign rv_inl24 = ((c1242 || c1243) || c1235) ? sub_add_result1_inl25 : ((c1250 || c1251) || c1244) ? sub_add_result2_inl25 : 'bz;
  assign rv_inl2_inl15 = ((c1262 || c1263) || c1259) ? sub_add_result1_inl2_inl16 : ((c1266 || c1267) || c1264) ? sub_add_result2_inl2_inl16 : 'bz;
  assign rv_n_inl1_inl22 = (t569_inl2 + t570_inl2);
  assign rv_n_inl1_inl23 = (rv_n_inl1_inl22 >>> 1);
  assign rv_n_inl1_inl24 = c1221 ? rv_n_inl1_inl23 : (c1216 && !c591_inl1_inl2) ? rv_n_inl1_inl22 : 'bz;
  assign rv_n_inl1_inl25 = (x_inl1_inl24 - b_inl1_inl24);
  assign rv_n_inl1_inl27 = (rv_n_inl1_inl26 << 1);
  assign rv_n_inl1_inl2_inl13 = (t569_inl2_inl1 + t570_inl2_inl1);
  assign rv_n_inl1_inl2_inl14 = (rv_n_inl1_inl2_inl13 >>> 1);
  assign rv_n_inl1_inl2_inl15 = c1246 ? rv_n_inl1_inl2_inl14 : (c1238 && !c591_inl1_inl2_inl1) ? rv_n_inl1_inl2_inl13 : 'bz;
  assign rv_n_inl1_inl2_inl16 = (x_inl1_inl2_inl15 - b_inl1_inl2_inl15);
  assign rv_n_inl1_inl2_inl18 = (rv_n_inl1_inl2_inl17 << 1);
  assign rv_n_inl2_inl22 = (t577_inl2 + new_b_n_inl2);
  assign rv_n_inl2_inl23 = (rv_n_inl2_inl22 >>> 1);
  assign rv_n_inl2_inl24 = c1227 ? rv_n_inl2_inl23 : (c1223 && !c591_inl2_inl2) ? rv_n_inl2_inl22 : 'bz;
  assign rv_n_inl2_inl25 = (x_inl2_inl24 - b_inl2_inl24);
  assign rv_n_inl2_inl27 = (rv_n_inl2_inl26 << 1);
  assign rv_n_inl2_inl2_inl13 = (t577_inl2_inl1 + new_b_n_inl2_inl1);
  assign rv_n_inl2_inl2_inl14 = (rv_n_inl2_inl2_inl13 >>> 1);
  assign rv_n_inl2_inl2_inl15 = c1253 ? rv_n_inl2_inl2_inl14 : (c1248 && !c591_inl2_inl2_inl1) ? rv_n_inl2_inl2_inl13 : 'bz;
  assign rv_n_inl2_inl2_inl16 = (x_inl2_inl2_inl15 - b_inl2_inl2_inl15);
  assign rv_n_inl2_inl2_inl18 = (rv_n_inl2_inl2_inl17 << 1);
  assign s_inl1_inl1 = (t626_inl1_inl1 ^ t627_inl1_inl1);
  assign sub_add_result1_inl22 = (t595_inl1_inl2 | t596_inl1_inl2);
  assign sub_add_result1_inl23 = (t603_inl1_inl2 | t604_inl1_inl2);
  assign sub_add_result1_inl25 = (c1226 || c1221) ? sub_add_result1_inl22 : c1235 ? sub_add_result1_inl23 : (c1222 || c1217) ? 0 : 'bz;
  assign sub_add_result1_inl2_inl13 = (t595_inl1_inl2_inl1 | t596_inl1_inl2_inl1);
  assign sub_add_result1_inl2_inl14 = (t603_inl1_inl2_inl1 | t604_inl1_inl2_inl1);
  assign sub_add_result1_inl2_inl16 = (c1252 || c1246) ? sub_add_result1_inl2_inl13 : c1259 ? sub_add_result1_inl2_inl14 : (c1247 || c1239) ? 0 : 'bz;
  assign sub_add_result2_inl22 = (t595_inl2_inl2 | t596_inl2_inl2);
  assign sub_add_result2_inl23 = (t603_inl2_inl2 | t604_inl2_inl2);
  assign sub_add_result2_inl25 = (c1232 || c1227) ? sub_add_result2_inl22 : c1244 ? sub_add_result2_inl23 : (c1228 || c1224) ? 0 : 'bz;
  assign sub_add_result2_inl2_inl13 = (t595_inl2_inl2_inl1 | t596_inl2_inl2_inl1);
  assign sub_add_result2_inl2_inl14 = (t603_inl2_inl2_inl1 | t604_inl2_inl2_inl1);
  assign sub_add_result2_inl2_inl16 = (c1258 || c1253) ? sub_add_result2_inl2_inl13 : c1264 ? sub_add_result2_inl2_inl14 : (c1254 || c1249) ? 0 : 'bz;
  assign t560_inl2 = (t612 & 32768);
  assign t560_inl2_inl1 = (mul_result1_inl16 & 32768);
  assign t561_inl2 = t560_inl2 ? 1 : 0;
  assign t561_inl2_inl1 = t560_inl2_inl1 ? 1 : 0;
  assign t562_inl2 = (t613 & 32768);
  assign t562_inl2_inl1 = (t609 & 32768);
  assign t563_inl2 = t562_inl2 ? 1 : 0;
  assign t563_inl2_inl1 = t562_inl2_inl1 ? 1 : 0;
  assign t564_inl2 = (t612 >>> 7);
  assign t564_inl2_inl1 = (mul_result1_inl16 >>> 7);
  assign t565_inl2 = (t613 >>> 7);
  assign t565_inl2_inl1 = (t609 >>> 7);
  assign t569_inl2 = (128 | x_n_inl2);
  assign t569_inl2_inl1 = (128 | x_n_inl2_inl1);
  assign t570_inl2 = (128 | b_n_inl2);
  assign t570_inl2_inl1 = (128 | b_n_inl2_inl1);
  assign t571_inl2 = (128 | b_n_inl2);
  assign t571_inl2_inl1 = (128 | b_n_inl2_inl1);
  assign t572_inl2 = (t571_inl2 >>> d_inl2);
  assign t572_inl2_inl1 = (t571_inl2_inl1 >>> d_inl2_inl1);
  assign t573_inl2 = (d_inl2 - 1);
  assign t573_inl2_inl1 = (d_inl2_inl1 - 1);
  assign t574_inl2 = (b_n_inl2 >>> t573_inl2);
  assign t574_inl2_inl1 = (b_n_inl2_inl1 >>> t573_inl2_inl1);
  assign t575_inl2 = (t574_inl2 & 1);
  assign t575_inl2_inl1 = (t574_inl2_inl1 & 1);
  assign t577_inl2 = (128 | x_n_inl2);
  assign t577_inl2_inl1 = (128 | x_n_inl2_inl1);
  assign t589_inl1_inl2 = (rv_n_inl1_inl22 & 256);
  assign t589_inl1_inl2_inl1 = (rv_n_inl1_inl2_inl13 & 256);
  assign t589_inl2_inl2 = (rv_n_inl2_inl22 & 256);
  assign t589_inl2_inl2_inl1 = (rv_n_inl2_inl2_inl13 & 256);
  assign t590_inl1_inl2 = t589_inl1_inl2 ? 1 : 0;
  assign t590_inl1_inl2_inl1 = t589_inl1_inl2_inl1 ? 1 : 0;
  assign t590_inl2_inl2 = t589_inl2_inl2 ? 1 : 0;
  assign t590_inl2_inl2_inl1 = t589_inl2_inl2_inl1 ? 1 : 0;
  assign t592_inl1_inl2 = x_sign_inl24 ? 32768 : 0;
  assign t592_inl1_inl2_inl1 = x_sign_inl2_inl15 ? 32768 : 0;
  assign t592_inl2_inl2 = x_sign_inl24 ? 32768 : 0;
  assign t592_inl2_inl2_inl1 = x_sign_inl2_inl15 ? 32768 : 0;
  assign t593_inl1_inl2 = (e_inl1_inl2 + t590_inl1_inl2);
  assign t593_inl1_inl2_inl1 = (e_inl1_inl2_inl1 + t590_inl1_inl2_inl1);
  assign t593_inl2_inl2 = (e_inl2_inl2 + t590_inl2_inl2);
  assign t593_inl2_inl2_inl1 = (e_inl2_inl2_inl1 + t590_inl2_inl2_inl1);
  assign t594_inl1_inl2 = (t593_inl1_inl2 << 7);
  assign t594_inl1_inl2_inl1 = (t593_inl1_inl2_inl1 << 7);
  assign t594_inl2_inl2 = (t593_inl2_inl2 << 7);
  assign t594_inl2_inl2_inl1 = (t593_inl2_inl2_inl1 << 7);
  assign t595_inl1_inl2 = (t592_inl1_inl2 | t594_inl1_inl2);
  assign t595_inl1_inl2_inl1 = (t592_inl1_inl2_inl1 | t594_inl1_inl2_inl1);
  assign t595_inl2_inl2 = (t592_inl2_inl2 | t594_inl2_inl2);
  assign t595_inl2_inl2_inl1 = (t592_inl2_inl2_inl1 | t594_inl2_inl2_inl1);
  assign t596_inl1_inl2 = (rv_n_inl1_inl24 & 127);
  assign t596_inl1_inl2_inl1 = (rv_n_inl1_inl2_inl15 & 127);
  assign t596_inl2_inl2 = (rv_n_inl2_inl24 & 127);
  assign t596_inl2_inl2_inl1 = (rv_n_inl2_inl2_inl15 & 127);
  assign t598_inl1_inl2 = (rv_n_inl1_inl26 & 128);
  assign t598_inl1_inl2_inl1 = (rv_n_inl1_inl2_inl17 & 128);
  assign t598_inl2_inl2 = (rv_n_inl2_inl26 & 128);
  assign t598_inl2_inl2_inl1 = (rv_n_inl2_inl2_inl17 & 128);
  assign t600_inl1_inl2 = x_sign_inl1_inl24 ? 32768 : 0;
  assign t600_inl1_inl2_inl1 = x_sign_inl1_inl2_inl15 ? 32768 : 0;
  assign t600_inl2_inl2 = x_sign_inl2_inl24 ? 32768 : 0;
  assign t600_inl2_inl2_inl1 = x_sign_inl2_inl2_inl15 ? 32768 : 0;
  assign t601_inl1_inl2 = (e_inl1_inl2 - i_inl1_inl23);
  assign t601_inl1_inl2_inl1 = (e_inl1_inl2_inl1 - i_inl1_inl2_inl14);
  assign t601_inl2_inl2 = (e_inl2_inl2 - i_inl2_inl23);
  assign t601_inl2_inl2_inl1 = (e_inl2_inl2_inl1 - i_inl2_inl2_inl14);
  assign t602_inl1_inl2 = (t601_inl1_inl2 << 7);
  assign t602_inl1_inl2_inl1 = (t601_inl1_inl2_inl1 << 7);
  assign t602_inl2_inl2 = (t601_inl2_inl2 << 7);
  assign t602_inl2_inl2_inl1 = (t601_inl2_inl2_inl1 << 7);
  assign t603_inl1_inl2 = (t600_inl1_inl2 | t602_inl1_inl2);
  assign t603_inl1_inl2_inl1 = (t600_inl1_inl2_inl1 | t602_inl1_inl2_inl1);
  assign t603_inl2_inl2 = (t600_inl2_inl2 | t602_inl2_inl2);
  assign t603_inl2_inl2_inl1 = (t600_inl2_inl2_inl1 | t602_inl2_inl2_inl1);
  assign t604_inl1_inl2 = (rv_n_inl1_inl26 & 127);
  assign t604_inl1_inl2_inl1 = (rv_n_inl1_inl2_inl17 & 127);
  assign t604_inl2_inl2 = (rv_n_inl2_inl26 & 127);
  assign t604_inl2_inl2_inl1 = (rv_n_inl2_inl2_inl17 & 127);
  assign t607 = (xi2 + j3);
  assign t608 = W_PARAM(t607);
  assign t613 = B_PARAM(j6);
  assign t617_inl1_inl1 = (x >>> 7);
  assign t618_inl1_inl1 = (t608 >>> 7);
  assign t619_inl1_inl1 = (x_e_inl1_inl1 - 127);
  assign t620_inl1_inl1 = (w_e_inl1_inl1 - 127);
  assign t621_inl1_inl1 = (t619_inl1_inl1 + t620_inl1_inl1);
  assign t622_inl1_inl1 = (x_n_inl1_inl1 | 128);
  assign t623_inl1_inl1 = (w_n_inl1_inl1 | 128);
  assign t624_inl1_inl1 = (new_n_inl1_inl13 & 32768);
  assign t626_inl1_inl1 = (x & 32768);
  assign t627_inl1_inl1 = (t608 & 32768);
  assign t628_inl1_inl1 = (e_inl1_inl15 << 7);
  assign t629_inl1_inl1 = (s_inl1_inl1 | t628_inl1_inl1);
  assign w_e_inl1_inl1 = (t618_inl1_inl1 & 255);
  assign w_n_inl1_inl1 = (t608 & 127);
  assign x_e_inl1_inl1 = (t617_inl1_inl1 & 255);
  assign x_e_inl22 = (t564_inl2 & 255);
  assign x_e_inl24 = c1206 ? b_e_inl22 : (c1203 && !c566_inl2) ? x_e_inl22 : 'bz;
  assign x_e_inl2_inl13 = (t564_inl2_inl1 & 255);
  assign x_e_inl2_inl15 = c1220 ? b_e_inl2_inl13 : (c1215 && !c566_inl2_inl1) ? x_e_inl2_inl13 : 'bz;
  assign x_inl1_inl24 = c1217 ? t570_inl2 : (c1212 && c644_inl1_inl2) ? t569_inl2 : 'bz;
  assign x_inl1_inl2_inl15 = c1239 ? t570_inl2_inl1 : (c1233 && c644_inl1_inl2_inl1) ? t569_inl2_inl1 : 'bz;
  assign x_inl24 = c1206 ? t613 : (c1203 && !c566_inl2) ? t612 : 'bz;
  assign x_inl2_inl15 = c1220 ? t609 : (c1215 && !c566_inl2_inl1) ? mul_result1_inl16 : 'bz;
  assign x_inl2_inl24 = c1224 ? new_b_n_inl2 : (c1219 && c644_inl2_inl2) ? t577_inl2 : 'bz;
  assign x_inl2_inl2_inl15 = c1249 ? new_b_n_inl2_inl1 : (c1241 && c644_inl2_inl2_inl1) ? t577_inl2_inl1 : 'bz;
  assign x_n_inl1_inl1 = (x & 127);
  assign x_n_inl2 = (x_inl24 & 127);
  assign x_n_inl2_inl1 = (x_inl2_inl15 & 127);
  assign x_sign_inl1_inl24 = c1217 ? b_sign_inl24 : (c1212 && c644_inl1_inl2) ? x_sign_inl24 : 'bz;
  assign x_sign_inl1_inl2_inl15 = c1239 ? b_sign_inl2_inl15 : (c1233 && c644_inl1_inl2_inl1) ? x_sign_inl2_inl15 : 'bz;
  assign x_sign_inl24 = c1206 ? t563_inl2 : (c1203 && !c566_inl2) ? t561_inl2 : 'bz;
  assign x_sign_inl2_inl15 = c1220 ? t563_inl2_inl1 : (c1215 && !c566_inl2_inl1) ? t561_inl2_inl1 : 'bz;
  assign x_sign_inl2_inl24 = c1224 ? b_sign_inl24 : (c1219 && c644_inl2_inl2) ? x_sign_inl24 : 'bz;
  assign x_sign_inl2_inl2_inl15 = c1249 ? b_sign_inl2_inl15 : (c1241 && c644_inl2_inl2_inl1) ? x_sign_inl2_inl15 : 'bz;
  assign x_w_inl1_inl1 = (t629_inl1_inl1 | new_n_inl1_inl17);
  assign xi3 = (xi2 + 10);
  //combinations: in__mem
  assign _mem_len = do_mnist7_mem_in__mem_len;
  assign _mem_q = do_mnist7_mem_in__mem_q;
  assign do_mnist7_mem_in__mem_addr = _mem_addr;
  assign do_mnist7_mem_in__mem_d = _mem_d;
  assign do_mnist7_mem_in__mem_req = _mem_req;
  assign do_mnist7_mem_in__mem_we = _mem_we;
  //combinations: in_a
  assign a_len = do_mnist7_mem_in_a_len;
  assign a_q = do_mnist7_mem_in_a_q;
  assign do_mnist7_mem_in_a_addr = a_addr;
  assign do_mnist7_mem_in_a_d = a_d;
  assign do_mnist7_mem_in_a_req = a_req;
  assign do_mnist7_mem_in_a_we = a_we;
  
  always @(posedge clk) begin
    if (rst) begin
      _mem_addr <= 0;
      _mem_d <= 0;
      _mem_req <= 0;
      _mem_we <= 0;
      a_addr <= 0;
      a_d <= 0;
      a_req <= 0;
      a_we <= 0;
      i2 <= 0;
      i_inl1_inl23 <= 0;
      i_inl1_inl2_inl14 <= 0;
      i_inl2_inl23 <= 0;
      i_inl2_inl2_inl14 <= 0;
      j3 <= 0;
      j6 <= 0;
      lst_len <= 0;
      rv_n_inl1_inl26 <= 0;
      rv_n_inl1_inl2_inl17 <= 0;
      rv_n_inl2_inl26 <= 0;
      rv_n_inl2_inl2_inl17 <= 0;
      t609 <= 0;
      t612 <= 0;
      x <= 0;
      xi2 <= 0;
      do_mnist7_mem_state <= do_mnist7_mem_b1_INIT;
    end else begin //if (rst)
      case(do_mnist7_mem_state)
      do_mnist7_mem_b1_INIT: begin
        do_mnist7_mem_valid <= 0;
        if (do_mnist7_mem_ready == 1) begin
          lst_len <= do_mnist7_mem_in_lst_len;
          array630[0] <= 0;
          array630[1] <= 0;
          array630[2] <= 0;
          array630[3] <= 0;
          array630[4] <= 0;
          array630[5] <= 0;
          array630[6] <= 0;
          array630[7] <= 0;
          array630[8] <= 0;
          array630[9] <= 0;
          i2 <= 0;
          xi2 <= 0;
          do_mnist7_mem_state <= do_mnist7_mem_L1_fortest2_S0;
        end
      end
      do_mnist7_mem_L1_fortest2_S0: begin
        /* c605 <= (i2 < lst_len); */
        j6 <= 0;
        do_mnist7_mem_state <= do_mnist7_mem_L1_fortest2_S1;
      end
      do_mnist7_mem_L1_fortest2_S1: begin
        if (c605) begin
          a_addr <= i2;
          a_we <= 0;
          a_req <= 1;
          j3 <= 0;
          do_mnist7_mem_state <= do_mnist7_mem_L1_forbody3_S1;
        end else begin
          /* c611 <= (j6 < 10); */
          if (c611) begin
            t612 <= array630[j6];
            /* t613 <= B_PARAM(j6); */
            do_mnist7_mem_state <= do_mnist7_mem_L5_forbody13_S1;
          end else begin
            do_mnist7_mem_valid <= 1;
            if (do_mnist7_mem_accept == 1) begin
              do_mnist7_mem_state <= do_mnist7_mem_b1_INIT;
            end
          end
        end
      end
      do_mnist7_mem_L1_forbody3_S1: begin
        /*wait for output of a*/
        do_mnist7_mem_state <= do_mnist7_mem_L1_forbody3_S2;
      end
      do_mnist7_mem_L1_forbody3_S2: begin
        x <= a_q;
        a_req <= 0;
        do_mnist7_mem_state <= do_mnist7_mem_L2_fortest4_S0;
      end
      do_mnist7_mem_L2_fortest4_S0: begin
        /* c606 <= (j3 < 10); */
        if (c606) begin
          /* t607 <= (xi2 + j3); */
          t609 <= array630[j3];
          /* c615_inl1_inl1 <= (x == 0); */
          /* t617_inl1_inl1 <= (x >>> 7); */
          /* x_n_inl1_inl1 <= (x & 127); */
          /* t626_inl1_inl1 <= (x & 32768); */
          /* c1677 <= (c605 && c606); */
          /* c1195 <= (c605 && c606); */
          /* t608 <= W_PARAM(t607); */
          /* x_e_inl1_inl1 <= (t617_inl1_inl1 & 255); */
          /* t622_inl1_inl1 <= (x_n_inl1_inl1 | 128); */
          /* c1196 <= (c1195 && c615_inl1_inl1); */
          /* c1197 <= (c1195 && !c615_inl1_inl1); */
          /* c616_inl1_inl1 <= (t608 == 0); */
          /* t618_inl1_inl1 <= (t608 >>> 7); */
          /* t619_inl1_inl1 <= (x_e_inl1_inl1 - 127); */
          /* w_n_inl1_inl1 <= (t608 & 127); */
          /* t627_inl1_inl1 <= (t608 & 32768); */
          /* c1200 <= (c1197 && c616_inl1_inl1); */
          /* c1201 <= (c1197 && !c616_inl1_inl1); */
          /* w_e_inl1_inl1 <= (t618_inl1_inl1 & 255); */
          /* t623_inl1_inl1 <= (w_n_inl1_inl1 | 128); */
          /* s_inl1_inl1 <= (t626_inl1_inl1 ^ t627_inl1_inl1); */
          /* t620_inl1_inl1 <= (w_e_inl1_inl1 - 127); */
          /* new_n_inl1_inl13 <= (t622_inl1_inl1 * t623_inl1_inl1); */
          /* t621_inl1_inl1 <= (t619_inl1_inl1 + t620_inl1_inl1); */
          /* t624_inl1_inl1 <= (new_n_inl1_inl13 & 32768); */
          /* new_n_inl1_inl14 <= (new_n_inl1_inl13 >>> 8); */
          /* new_n_inl1_inl15 <= (new_n_inl1_inl13 >>> 7); */
          /* e_inl1_inl13 <= (t621_inl1_inl1 + 127); */
          /* c625_inl1_inl1 <= (t624_inl1_inl1 != 0); */
          /* c1204 <= (c1201 && c625_inl1_inl1); */
          /* e_inl1_inl14 <= (e_inl1_inl13 + 1); */
          /* c1205 <= (c1201 && !c625_inl1_inl1); */
          /* e_inl1_inl15 <= c1204 ? e_inl1_inl14 : c1205 ? e_inl1_inl13 : 'bz; */
          /* new_n_inl1_inl16 <= c1204 ? new_n_inl1_inl14 : c1205 ? new_n_inl1_inl15 : 'bz; */
          /* new_n_inl1_inl17 <= (new_n_inl1_inl16 & 127); */
          /* t628_inl1_inl1 <= (e_inl1_inl15 << 7); */
          /* t629_inl1_inl1 <= (s_inl1_inl1 | t628_inl1_inl1); */
          /* x_w_inl1_inl1 <= (t629_inl1_inl1 | new_n_inl1_inl17); */
          /* mul_result1_inl16 <= c1196 ? 0 : (c1197 && c1200) ? 0 : (c1197 && (c1205 || c1204)) ? x_w_inl1_inl1 : 'bz; */
          /* c558_inl2_inl1 <= (mul_result1_inl16 == 0); */
          new_n_inl1_inl13 <= (t622_inl1_inl1 * t623_inl1_inl1);
          do_mnist7_mem_state <= do_mnist7_mem_L2_forbody5_S1_MUL;
        end else begin
          /* xi3 <= (xi2 + 10); */
          /* i3 <= (i2 + 1); */
          i2 <= i3;
          xi2 <= xi3;
          do_mnist7_mem_state <= do_mnist7_mem_L1_fortest2_S0;
        end
      end
      do_mnist7_mem_L2_forbody5_S1_MUL: begin
        do_mnist7_mem_state <= do_mnist7_mem_L2_forbody5_S1;
      end
      do_mnist7_mem_L2_forbody5_S1: begin
        if (c558_inl2_inl1) begin
          /* c1680 <= (c1677 && c558_inl2_inl1); */
          /* c1210 <= (c1195 && c558_inl2_inl1); */
          do_mnist7_mem_state <= do_mnist7_mem_L2_exit25_S0;
        end else begin
          /* c559_inl2_inl1 <= (t609 == 0); */
          /* c1681 <= (c1677 && !c558_inl2_inl1); */
          /* c1211 <= (c1195 && !c558_inl2_inl1); */
          if (c559_inl2_inl1) begin
            /* c1684 <= (c1681 && c559_inl2_inl1); */
            /* c1214 <= (c1211 && c559_inl2_inl1); */
            do_mnist7_mem_state <= do_mnist7_mem_L2_exit25_S0;
          end else begin
            /* t562_inl2_inl1 <= (t609 & 32768); */
            /* t565_inl2_inl1 <= (t609 >>> 7); */
            /* t563_inl2_inl1 <= t562_inl2_inl1 ? 1 : 0; */
            /* b_e_inl2_inl13 <= (t565_inl2_inl1 & 255); */
            /* t560_inl2_inl1 <= (mul_result1_inl16 & 32768); */
            /* t564_inl2_inl1 <= (mul_result1_inl16 >>> 7); */
            /* t561_inl2_inl1 <= t560_inl2_inl1 ? 1 : 0; */
            /* x_e_inl2_inl13 <= (t564_inl2_inl1 & 255); */
            /* c1685 <= (c1681 && !c559_inl2_inl1); */
            /* c1215 <= (c1211 && !c559_inl2_inl1); */
            /* c566_inl2_inl1 <= (x_e_inl2_inl13 < b_e_inl2_inl13); */
            /* c1220 <= (c1215 && c566_inl2_inl1); */
            /* c1225 <= (c1215 && !c566_inl2_inl1); */
            /* b_e_inl2_inl15 <= c1220 ? x_e_inl2_inl13 : (c1215 && !c566_inl2_inl1) ? b_e_inl2_inl13 : 'bz; */
            /* b_inl2_inl15 <= c1220 ? mul_result1_inl16 : (c1215 && !c566_inl2_inl1) ? t609 : 'bz; */
            /* b_sign_inl2_inl15 <= c1220 ? t561_inl2_inl1 : (c1215 && !c566_inl2_inl1) ? t563_inl2_inl1 : 'bz; */
            /* x_e_inl2_inl15 <= c1220 ? b_e_inl2_inl13 : (c1215 && !c566_inl2_inl1) ? x_e_inl2_inl13 : 'bz; */
            /* x_inl2_inl15 <= c1220 ? t609 : (c1215 && !c566_inl2_inl1) ? mul_result1_inl16 : 'bz; */
            /* x_sign_inl2_inl15 <= c1220 ? t563_inl2_inl1 : (c1215 && !c566_inl2_inl1) ? t561_inl2_inl1 : 'bz; */
            /* x_n_inl2_inl1 <= (x_inl2_inl15 & 127); */
            /* b_n_inl2_inl1 <= (b_inl2_inl15 & 127); */
            /* d_inl2_inl1 <= (x_e_inl2_inl15 - b_e_inl2_inl15); */
            /* c567_inl2_inl1 <= (d_inl2_inl1 > 8); */
            if (c567_inl2_inl1) begin
              /* c1688 <= (c1685 && c567_inl2_inl1); */
              /* c1229 <= ((c1225 || c1220) && c567_inl2_inl1); */
              do_mnist7_mem_state <= do_mnist7_mem_L2_exit25_S0;
            end else begin
              /* c568_inl2_inl1 <= (d_inl2_inl1 == 0); */
              /* c1689 <= (c1685 && !c567_inl2_inl1); */
              /* c1230 <= ((c1225 || c1220) && !c567_inl2_inl1); */
              if (c568_inl2_inl1) begin
                /* e_inl1_inl2_inl1 <= x_e_inl2_inl15; */
                /* c581_inl1_inl2_inl1 <= (x_sign_inl2_inl15 == 0); */
                /* c582_inl1_inl2_inl1 <= (b_sign_inl2_inl15 == 0); */
                /* c584_inl1_inl2_inl1 <= (x_sign_inl2_inl15 == 1); */
                /* c585_inl1_inl2_inl1 <= (b_sign_inl2_inl15 == 1); */
                /* t569_inl2_inl1 <= (128 | x_n_inl2_inl1); */
                /* t570_inl2_inl1 <= (128 | b_n_inl2_inl1); */
                /* c583_inl1_inl2_inl1 <= (c581_inl1_inl2_inl1 && c582_inl1_inl2_inl1); */
                /* c586_inl1_inl2_inl1 <= (c584_inl1_inl2_inl1 && c585_inl1_inl2_inl1); */
                /* c587_inl1_inl2_inl1 <= (c583_inl1_inl2_inl1 || c586_inl1_inl2_inl1); */
                /* c588_inl1_inl2_inl1 <= (t569_inl2_inl1 < t570_inl2_inl1); */
                /* c1692 <= (c1689 && c568_inl2_inl1); */
                /* c1233 <= (c1230 && c568_inl2_inl1); */
                /* c643_inl1_inl2_inl1 <= (!c587_inl1_inl2_inl1 && c588_inl1_inl2_inl1); */
                /* c644_inl1_inl2_inl1 <= (!c587_inl1_inl2_inl1 && !c588_inl1_inl2_inl1); */
                if (c587_inl1_inl2_inl1) begin
                  /* t592_inl1_inl2_inl1 <= x_sign_inl2_inl15 ? 32768 : 0; */
                  /* rv_n_inl1_inl2_inl13 <= (t569_inl2_inl1 + t570_inl2_inl1); */
                  /* t589_inl1_inl2_inl1 <= (rv_n_inl1_inl2_inl13 & 256); */
                  /* rv_n_inl1_inl2_inl14 <= (rv_n_inl1_inl2_inl13 >>> 1); */
                  /* c1698 <= (c1692 && c587_inl1_inl2_inl1); */
                  /* c1238 <= (c1233 && c587_inl1_inl2_inl1); */
                  /* t590_inl1_inl2_inl1 <= t589_inl1_inl2_inl1 ? 1 : 0; */
                  /* c591_inl1_inl2_inl1 <= (t590_inl1_inl2_inl1 != 0); */
                  /* t593_inl1_inl2_inl1 <= (e_inl1_inl2_inl1 + t590_inl1_inl2_inl1); */
                  /* c1246 <= (c1238 && c591_inl1_inl2_inl1); */
                  /* c1252 <= (c1238 && !c591_inl1_inl2_inl1); */
                  /* t594_inl1_inl2_inl1 <= (t593_inl1_inl2_inl1 << 7); */
                  /* rv_n_inl1_inl2_inl15 <= c1246 ? rv_n_inl1_inl2_inl14 : (c1238 && !c591_inl1_inl2_inl1) ? rv_n_inl1_inl2_inl13 : 'bz; */
                  /* t595_inl1_inl2_inl1 <= (t592_inl1_inl2_inl1 | t594_inl1_inl2_inl1); */
                  /* t596_inl1_inl2_inl1 <= (rv_n_inl1_inl2_inl15 & 127); */
                  /* sub_add_result1_inl2_inl13 <= (t595_inl1_inl2_inl1 | t596_inl1_inl2_inl1); */
                  do_mnist7_mem_state <= do_mnist7_mem_L2_exit39_S0;
                end else begin
                  /* c1699 <= (c1692 && !c587_inl1_inl2_inl1); */
                  /* c1239 <= (c1233 && c643_inl1_inl2_inl1); */
                  do_mnist7_mem_state <= do_mnist7_mem_L2_b43_S0;
                end
              end else begin
                /* t571_inl2_inl1 <= (128 | b_n_inl2_inl1); */
                /* t573_inl2_inl1 <= (d_inl2_inl1 - 1); */
                /* t572_inl2_inl1 <= (t571_inl2_inl1 >>> d_inl2_inl1); */
                /* t574_inl2_inl1 <= (b_n_inl2_inl1 >>> t573_inl2_inl1); */
                /* c1693 <= (c1689 && !c568_inl2_inl1); */
                /* c1234 <= (c1230 && !c568_inl2_inl1); */
                /* t575_inl2_inl1 <= (t574_inl2_inl1 & 1); */
                /* new_b_n_inl2_inl1 <= (t572_inl2_inl1 + t575_inl2_inl1); */
                /* c576_inl2_inl1 <= (new_b_n_inl2_inl1 == 0); */
                if (c576_inl2_inl1) begin
                  /* c1700 <= (c1693 && c576_inl2_inl1); */
                  /* c1240 <= (c1234 && c576_inl2_inl1); */
                  do_mnist7_mem_state <= do_mnist7_mem_L2_exit25_S0;
                end else begin
                  /* e_inl2_inl2_inl1 <= x_e_inl2_inl15; */
                  /* c581_inl2_inl2_inl1 <= (x_sign_inl2_inl15 == 0); */
                  /* c582_inl2_inl2_inl1 <= (b_sign_inl2_inl15 == 0); */
                  /* c584_inl2_inl2_inl1 <= (x_sign_inl2_inl15 == 1); */
                  /* c585_inl2_inl2_inl1 <= (b_sign_inl2_inl15 == 1); */
                  /* t577_inl2_inl1 <= (128 | x_n_inl2_inl1); */
                  /* c583_inl2_inl2_inl1 <= (c581_inl2_inl2_inl1 && c582_inl2_inl2_inl1); */
                  /* c586_inl2_inl2_inl1 <= (c584_inl2_inl2_inl1 && c585_inl2_inl2_inl1); */
                  /* c587_inl2_inl2_inl1 <= (c583_inl2_inl2_inl1 || c586_inl2_inl2_inl1); */
                  /* c588_inl2_inl2_inl1 <= (t577_inl2_inl1 < new_b_n_inl2_inl1); */
                  /* c1701 <= (c1693 && !c576_inl2_inl1); */
                  /* c1241 <= (c1234 && !c576_inl2_inl1); */
                  /* c643_inl2_inl2_inl1 <= (!c587_inl2_inl2_inl1 && c588_inl2_inl2_inl1); */
                  /* c644_inl2_inl2_inl1 <= (!c587_inl2_inl2_inl1 && !c588_inl2_inl2_inl1); */
                  if (c587_inl2_inl2_inl1) begin
                    /* t592_inl2_inl2_inl1 <= x_sign_inl2_inl15 ? 32768 : 0; */
                    /* rv_n_inl2_inl2_inl13 <= (t577_inl2_inl1 + new_b_n_inl2_inl1); */
                    /* t589_inl2_inl2_inl1 <= (rv_n_inl2_inl2_inl13 & 256); */
                    /* rv_n_inl2_inl2_inl14 <= (rv_n_inl2_inl2_inl13 >>> 1); */
                    /* c1704 <= (c1701 && c587_inl2_inl2_inl1); */
                    /* c1248 <= (c1241 && c587_inl2_inl2_inl1); */
                    /* t590_inl2_inl2_inl1 <= t589_inl2_inl2_inl1 ? 1 : 0; */
                    /* c591_inl2_inl2_inl1 <= (t590_inl2_inl2_inl1 != 0); */
                    /* t593_inl2_inl2_inl1 <= (e_inl2_inl2_inl1 + t590_inl2_inl2_inl1); */
                    /* c1253 <= (c1248 && c591_inl2_inl2_inl1); */
                    /* c1258 <= (c1248 && !c591_inl2_inl2_inl1); */
                    /* t594_inl2_inl2_inl1 <= (t593_inl2_inl2_inl1 << 7); */
                    /* rv_n_inl2_inl2_inl15 <= c1253 ? rv_n_inl2_inl2_inl14 : (c1248 && !c591_inl2_inl2_inl1) ? rv_n_inl2_inl2_inl13 : 'bz; */
                    /* t595_inl2_inl2_inl1 <= (t592_inl2_inl2_inl1 | t594_inl2_inl2_inl1); */
                    /* t596_inl2_inl2_inl1 <= (rv_n_inl2_inl2_inl15 & 127); */
                    /* sub_add_result2_inl2_inl13 <= (t595_inl2_inl2_inl1 | t596_inl2_inl2_inl1); */
                    do_mnist7_mem_state <= do_mnist7_mem_L2_exit56_S0;
                  end else begin
                    /* c1705 <= (c1701 && !c587_inl2_inl2_inl1); */
                    /* c1249 <= (c1241 && c643_inl2_inl2_inl1); */
                    do_mnist7_mem_state <= do_mnist7_mem_L2_b59_S0;
                  end
                end
              end
            end
          end
        end
      end
      do_mnist7_mem_L2_b43_S0: begin
        i_inl1_inl2_inl14 <= 0;
        /* c1247 <= (c1233 && c644_inl1_inl2_inl1); */
        /* b_inl1_inl2_inl15 <= c1239 ? t569_inl2_inl1 : (c1233 && c644_inl1_inl2_inl1) ? t570_inl2_inl1 : 'bz; */
        /* x_inl1_inl2_inl15 <= c1239 ? t570_inl2_inl1 : (c1233 && c644_inl1_inl2_inl1) ? t569_inl2_inl1 : 'bz; */
        /* x_sign_inl1_inl2_inl15 <= c1239 ? b_sign_inl2_inl15 : (c1233 && c644_inl1_inl2_inl1) ? x_sign_inl2_inl15 : 'bz; */
        /* rv_n_inl1_inl2_inl16 <= (x_inl1_inl2_inl15 - b_inl1_inl2_inl15); */
        rv_n_inl1_inl2_inl17 <= rv_n_inl1_inl2_inl16;
        do_mnist7_mem_state <= do_mnist7_mem_L4_fortest44_S0;
      end
      do_mnist7_mem_L2_b59_S0: begin
        i_inl2_inl2_inl14 <= 0;
        /* c1254 <= (c1241 && c644_inl2_inl2_inl1); */
        /* b_inl2_inl2_inl15 <= c1249 ? t577_inl2_inl1 : (c1241 && c644_inl2_inl2_inl1) ? new_b_n_inl2_inl1 : 'bz; */
        /* x_inl2_inl2_inl15 <= c1249 ? new_b_n_inl2_inl1 : (c1241 && c644_inl2_inl2_inl1) ? t577_inl2_inl1 : 'bz; */
        /* x_sign_inl2_inl2_inl15 <= c1249 ? b_sign_inl2_inl15 : (c1241 && c644_inl2_inl2_inl1) ? x_sign_inl2_inl15 : 'bz; */
        /* rv_n_inl2_inl2_inl16 <= (x_inl2_inl2_inl15 - b_inl2_inl2_inl15); */
        rv_n_inl2_inl2_inl17 <= rv_n_inl2_inl2_inl16;
        do_mnist7_mem_state <= do_mnist7_mem_L3_fortest60_S0;
      end
      do_mnist7_mem_L2_exit39_S0: begin
        /* c1717 <= (c1699 && !c597_inl1_inl2_inl1); */
        /* c1263 <= (c1247 || c1239); */
        /* c1262 <= (c1252 || c1246); */
        /* sub_add_result1_inl2_inl16 <= (c1252 || c1246) ? sub_add_result1_inl2_inl13 : c1259 ? sub_add_result1_inl2_inl14 : (c1247 || c1239) ? 0 : 'bz; */
        do_mnist7_mem_state <= do_mnist7_mem_L2_b41_S0;
      end
      do_mnist7_mem_L2_exit56_S0: begin
        /* c1721 <= (c1705 && !c597_inl2_inl2_inl1); */
        /* c1267 <= (c1254 || c1249); */
        /* c1266 <= (c1258 || c1253); */
        /* sub_add_result2_inl2_inl16 <= (c1258 || c1253) ? sub_add_result2_inl2_inl13 : c1264 ? sub_add_result2_inl2_inl14 : (c1254 || c1249) ? 0 : 'bz; */
        do_mnist7_mem_state <= do_mnist7_mem_L2_b41_S0;
      end
      do_mnist7_mem_L2_b41_S0: begin
        /* c1724 <= ((c1698 || c1717) || c1711); */
        /* c1268 <= ((c1262 || c1263) || c1259); */
        /* c1725 <= ((c1704 || c1721) || c1718); */
        /* c1269 <= ((c1266 || c1267) || c1264); */
        /* rv_inl2_inl15 <= ((c1262 || c1263) || c1259) ? sub_add_result1_inl2_inl16 : ((c1266 || c1267) || c1264) ? sub_add_result2_inl2_inl16 : 'bz; */
        /* add_result2_inl17 <= rv_inl2_inl15; */
        do_mnist7_mem_state <= do_mnist7_mem_L2_exit25_S0;
      end
      do_mnist7_mem_L2_exit25_S0: begin
        /* j4 <= (j3 + 1); */
        /* add_result2_inl18 <= c1210 ? t609 : c1214 ? mul_result1_inl16 : c1229 ? x_inl2_inl15 : c1240 ? x_inl2_inl15 : (c1268 || c1269) ? add_result2_inl17 : 'bz; */
        array630[j3] <= add_result2_inl18;
        j3 <= j4;
        do_mnist7_mem_state <= do_mnist7_mem_L2_fortest4_S0;
      end
      do_mnist7_mem_L3_fortest60_S0: begin
        /* c597_inl2_inl2_inl1 <= (i_inl2_inl2_inl14 < 7); */
        if (c597_inl2_inl2_inl1) begin
          /* t598_inl2_inl2_inl1 <= (rv_n_inl2_inl2_inl17 & 128); */
          /* c1713 <= (c1705 && c597_inl2_inl2_inl1); */
          /* c1261 <= ((c1254 || c1249) && c597_inl2_inl2_inl1); */
          /* c599_inl2_inl2_inl1 <= (t598_inl2_inl2_inl1 != 0); */
          if (c599_inl2_inl2_inl1) begin
            /* c1718 <= (c1713 && c599_inl2_inl2_inl1); */
            /* c1264 <= (c1261 && c599_inl2_inl2_inl1); */
            /* t601_inl2_inl2_inl1 <= (e_inl2_inl2_inl1 - i_inl2_inl2_inl14); */
            /* t602_inl2_inl2_inl1 <= (t601_inl2_inl2_inl1 << 7); */
            /* t600_inl2_inl2_inl1 <= x_sign_inl2_inl2_inl15 ? 32768 : 0; */
            /* t603_inl2_inl2_inl1 <= (t600_inl2_inl2_inl1 | t602_inl2_inl2_inl1); */
            /* t604_inl2_inl2_inl1 <= (rv_n_inl2_inl2_inl17 & 127); */
            /* sub_add_result2_inl2_inl14 <= (t603_inl2_inl2_inl1 | t604_inl2_inl2_inl1); */
            do_mnist7_mem_state <= do_mnist7_mem_L2_exit56_S0;
          end else begin
            /* rv_n_inl2_inl2_inl18 <= (rv_n_inl2_inl2_inl17 << 1); */
            /* i_inl2_inl2_inl15 <= (i_inl2_inl2_inl14 + 1); */
            i_inl2_inl2_inl14 <= i_inl2_inl2_inl15;
            rv_n_inl2_inl2_inl17 <= rv_n_inl2_inl2_inl18;
            /* c1719 <= (c1713 && !c599_inl2_inl2_inl1); */
            /* c1265 <= (c1261 && !c599_inl2_inl2_inl1); */
            do_mnist7_mem_state <= do_mnist7_mem_L3_fortest60_S0;
          end
        end else begin
          /* c1721 <= (c1705 && !c597_inl2_inl2_inl1); */
          /* c1267 <= (c1254 || c1249); */
          /* c1266 <= (c1258 || c1253); */
          /* sub_add_result2_inl2_inl16 <= (c1258 || c1253) ? sub_add_result2_inl2_inl13 : c1264 ? sub_add_result2_inl2_inl14 : (c1254 || c1249) ? 0 : 'bz; */
          do_mnist7_mem_state <= do_mnist7_mem_L2_b41_S0;
        end
      end
      do_mnist7_mem_L4_fortest44_S0: begin
        /* c597_inl1_inl2_inl1 <= (i_inl1_inl2_inl14 < 7); */
        if (c597_inl1_inl2_inl1) begin
          /* t598_inl1_inl2_inl1 <= (rv_n_inl1_inl2_inl17 & 128); */
          /* c1707 <= (c1699 && c597_inl1_inl2_inl1); */
          /* c1257 <= ((c1247 || c1239) && c597_inl1_inl2_inl1); */
          /* c599_inl1_inl2_inl1 <= (t598_inl1_inl2_inl1 != 0); */
          if (c599_inl1_inl2_inl1) begin
            /* c1711 <= (c1707 && c599_inl1_inl2_inl1); */
            /* c1259 <= (c1257 && c599_inl1_inl2_inl1); */
            /* t601_inl1_inl2_inl1 <= (e_inl1_inl2_inl1 - i_inl1_inl2_inl14); */
            /* t602_inl1_inl2_inl1 <= (t601_inl1_inl2_inl1 << 7); */
            /* t600_inl1_inl2_inl1 <= x_sign_inl1_inl2_inl15 ? 32768 : 0; */
            /* t603_inl1_inl2_inl1 <= (t600_inl1_inl2_inl1 | t602_inl1_inl2_inl1); */
            /* t604_inl1_inl2_inl1 <= (rv_n_inl1_inl2_inl17 & 127); */
            /* sub_add_result1_inl2_inl14 <= (t603_inl1_inl2_inl1 | t604_inl1_inl2_inl1); */
            do_mnist7_mem_state <= do_mnist7_mem_L2_exit39_S0;
          end else begin
            /* rv_n_inl1_inl2_inl18 <= (rv_n_inl1_inl2_inl17 << 1); */
            /* i_inl1_inl2_inl15 <= (i_inl1_inl2_inl14 + 1); */
            i_inl1_inl2_inl14 <= i_inl1_inl2_inl15;
            rv_n_inl1_inl2_inl17 <= rv_n_inl1_inl2_inl18;
            /* c1712 <= (c1707 && !c599_inl1_inl2_inl1); */
            /* c1260 <= (c1257 && !c599_inl1_inl2_inl1); */
            do_mnist7_mem_state <= do_mnist7_mem_L4_fortest44_S0;
          end
        end else begin
          /* c1717 <= (c1699 && !c597_inl1_inl2_inl1); */
          /* c1263 <= (c1247 || c1239); */
          /* c1262 <= (c1252 || c1246); */
          /* sub_add_result1_inl2_inl16 <= (c1252 || c1246) ? sub_add_result1_inl2_inl13 : c1259 ? sub_add_result1_inl2_inl14 : (c1247 || c1239) ? 0 : 'bz; */
          do_mnist7_mem_state <= do_mnist7_mem_L2_b41_S0;
        end
      end
      do_mnist7_mem_L5_fortest12_S0: begin
        /* c611 <= (j6 < 10); */
        if (c611) begin
          t612 <= array630[j6];
          /* t613 <= B_PARAM(j6); */
          do_mnist7_mem_state <= do_mnist7_mem_L5_forbody13_S1;
        end else begin
          do_mnist7_mem_valid <= 1;
          if (do_mnist7_mem_accept == 1) begin
            do_mnist7_mem_state <= do_mnist7_mem_b1_INIT;
          end
        end
      end
      do_mnist7_mem_L5_forbody13_S1: begin
        /* c558_inl2 <= (t612 == 0); */
        if (c558_inl2) begin
          /* c1678 <= (c611 && c558_inl2); */
          /* c1198 <= (c611 && c558_inl2); */
          do_mnist7_mem_state <= do_mnist7_mem_L5_exit74_S0;
        end else begin
          /* c559_inl2 <= (t613 == 0); */
          /* c1679 <= (c611 && !c558_inl2); */
          /* c1199 <= (c611 && !c558_inl2); */
          if (c559_inl2) begin
            /* c1682 <= (c1679 && c559_inl2); */
            /* c1202 <= (c1199 && c559_inl2); */
            do_mnist7_mem_state <= do_mnist7_mem_L5_exit74_S0;
          end else begin
            /* t560_inl2 <= (t612 & 32768); */
            /* t562_inl2 <= (t613 & 32768); */
            /* t564_inl2 <= (t612 >>> 7); */
            /* t565_inl2 <= (t613 >>> 7); */
            /* t561_inl2 <= t560_inl2 ? 1 : 0; */
            /* t563_inl2 <= t562_inl2 ? 1 : 0; */
            /* x_e_inl22 <= (t564_inl2 & 255); */
            /* b_e_inl22 <= (t565_inl2 & 255); */
            /* c1683 <= (c1679 && !c559_inl2); */
            /* c1203 <= (c1199 && !c559_inl2); */
            /* c566_inl2 <= (x_e_inl22 < b_e_inl22); */
            /* c1206 <= (c1203 && c566_inl2); */
            /* c1207 <= (c1203 && !c566_inl2); */
            /* b_e_inl24 <= c1206 ? x_e_inl22 : (c1203 && !c566_inl2) ? b_e_inl22 : 'bz; */
            /* b_inl24 <= c1206 ? t612 : (c1203 && !c566_inl2) ? t613 : 'bz; */
            /* b_sign_inl24 <= c1206 ? t561_inl2 : (c1203 && !c566_inl2) ? t563_inl2 : 'bz; */
            /* x_e_inl24 <= c1206 ? b_e_inl22 : (c1203 && !c566_inl2) ? x_e_inl22 : 'bz; */
            /* x_inl24 <= c1206 ? t613 : (c1203 && !c566_inl2) ? t612 : 'bz; */
            /* x_sign_inl24 <= c1206 ? t563_inl2 : (c1203 && !c566_inl2) ? t561_inl2 : 'bz; */
            /* x_n_inl2 <= (x_inl24 & 127); */
            /* b_n_inl2 <= (b_inl24 & 127); */
            /* d_inl2 <= (x_e_inl24 - b_e_inl24); */
            /* c567_inl2 <= (d_inl2 > 8); */
            if (c567_inl2) begin
              /* c1686 <= (c1683 && c567_inl2); */
              /* c1208 <= ((c1207 || c1206) && c567_inl2); */
              do_mnist7_mem_state <= do_mnist7_mem_L5_exit74_S0;
            end else begin
              /* c568_inl2 <= (d_inl2 == 0); */
              /* c1687 <= (c1683 && !c567_inl2); */
              /* c1209 <= ((c1207 || c1206) && !c567_inl2); */
              if (c568_inl2) begin
                /* e_inl1_inl2 <= x_e_inl24; */
                /* c581_inl1_inl2 <= (x_sign_inl24 == 0); */
                /* c582_inl1_inl2 <= (b_sign_inl24 == 0); */
                /* c584_inl1_inl2 <= (x_sign_inl24 == 1); */
                /* c585_inl1_inl2 <= (b_sign_inl24 == 1); */
                /* t569_inl2 <= (128 | x_n_inl2); */
                /* t570_inl2 <= (128 | b_n_inl2); */
                /* c583_inl1_inl2 <= (c581_inl1_inl2 && c582_inl1_inl2); */
                /* c586_inl1_inl2 <= (c584_inl1_inl2 && c585_inl1_inl2); */
                /* c587_inl1_inl2 <= (c583_inl1_inl2 || c586_inl1_inl2); */
                /* c588_inl1_inl2 <= (t569_inl2 < t570_inl2); */
                /* c1690 <= (c1687 && c568_inl2); */
                /* c1212 <= (c1209 && c568_inl2); */
                /* c643_inl1_inl2 <= (!c587_inl1_inl2 && c588_inl1_inl2); */
                /* c644_inl1_inl2 <= (!c587_inl1_inl2 && !c588_inl1_inl2); */
                if (c587_inl1_inl2) begin
                  /* t592_inl1_inl2 <= x_sign_inl24 ? 32768 : 0; */
                  /* rv_n_inl1_inl22 <= (t569_inl2 + t570_inl2); */
                  /* t589_inl1_inl2 <= (rv_n_inl1_inl22 & 256); */
                  /* rv_n_inl1_inl23 <= (rv_n_inl1_inl22 >>> 1); */
                  /* c1694 <= (c1690 && c587_inl1_inl2); */
                  /* c1216 <= (c1212 && c587_inl1_inl2); */
                  /* t590_inl1_inl2 <= t589_inl1_inl2 ? 1 : 0; */
                  /* c591_inl1_inl2 <= (t590_inl1_inl2 != 0); */
                  /* t593_inl1_inl2 <= (e_inl1_inl2 + t590_inl1_inl2); */
                  /* c1221 <= (c1216 && c591_inl1_inl2); */
                  /* c1226 <= (c1216 && !c591_inl1_inl2); */
                  /* t594_inl1_inl2 <= (t593_inl1_inl2 << 7); */
                  /* rv_n_inl1_inl24 <= c1221 ? rv_n_inl1_inl23 : (c1216 && !c591_inl1_inl2) ? rv_n_inl1_inl22 : 'bz; */
                  /* t595_inl1_inl2 <= (t592_inl1_inl2 | t594_inl1_inl2); */
                  /* t596_inl1_inl2 <= (rv_n_inl1_inl24 & 127); */
                  /* sub_add_result1_inl22 <= (t595_inl1_inl2 | t596_inl1_inl2); */
                  do_mnist7_mem_state <= do_mnist7_mem_L5_exit87_S0;
                end else begin
                  /* c1695 <= (c1690 && !c587_inl1_inl2); */
                  /* c1217 <= (c1212 && c643_inl1_inl2); */
                  do_mnist7_mem_state <= do_mnist7_mem_L5_b91_S0;
                end
              end else begin
                /* t571_inl2 <= (128 | b_n_inl2); */
                /* t573_inl2 <= (d_inl2 - 1); */
                /* t572_inl2 <= (t571_inl2 >>> d_inl2); */
                /* t574_inl2 <= (b_n_inl2 >>> t573_inl2); */
                /* c1691 <= (c1687 && !c568_inl2); */
                /* c1213 <= (c1209 && !c568_inl2); */
                /* t575_inl2 <= (t574_inl2 & 1); */
                /* new_b_n_inl2 <= (t572_inl2 + t575_inl2); */
                /* c576_inl2 <= (new_b_n_inl2 == 0); */
                if (c576_inl2) begin
                  /* c1696 <= (c1691 && c576_inl2); */
                  /* c1218 <= (c1213 && c576_inl2); */
                  do_mnist7_mem_state <= do_mnist7_mem_L5_exit74_S0;
                end else begin
                  /* e_inl2_inl2 <= x_e_inl24; */
                  /* c581_inl2_inl2 <= (x_sign_inl24 == 0); */
                  /* c582_inl2_inl2 <= (b_sign_inl24 == 0); */
                  /* c584_inl2_inl2 <= (x_sign_inl24 == 1); */
                  /* c585_inl2_inl2 <= (b_sign_inl24 == 1); */
                  /* t577_inl2 <= (128 | x_n_inl2); */
                  /* c583_inl2_inl2 <= (c581_inl2_inl2 && c582_inl2_inl2); */
                  /* c586_inl2_inl2 <= (c584_inl2_inl2 && c585_inl2_inl2); */
                  /* c587_inl2_inl2 <= (c583_inl2_inl2 || c586_inl2_inl2); */
                  /* c588_inl2_inl2 <= (t577_inl2 < new_b_n_inl2); */
                  /* c1697 <= (c1691 && !c576_inl2); */
                  /* c1219 <= (c1213 && !c576_inl2); */
                  /* c643_inl2_inl2 <= (!c587_inl2_inl2 && c588_inl2_inl2); */
                  /* c644_inl2_inl2 <= (!c587_inl2_inl2 && !c588_inl2_inl2); */
                  if (c587_inl2_inl2) begin
                    /* t592_inl2_inl2 <= x_sign_inl24 ? 32768 : 0; */
                    /* rv_n_inl2_inl22 <= (t577_inl2 + new_b_n_inl2); */
                    /* t589_inl2_inl2 <= (rv_n_inl2_inl22 & 256); */
                    /* rv_n_inl2_inl23 <= (rv_n_inl2_inl22 >>> 1); */
                    /* c1702 <= (c1697 && c587_inl2_inl2); */
                    /* c1223 <= (c1219 && c587_inl2_inl2); */
                    /* t590_inl2_inl2 <= t589_inl2_inl2 ? 1 : 0; */
                    /* c591_inl2_inl2 <= (t590_inl2_inl2 != 0); */
                    /* t593_inl2_inl2 <= (e_inl2_inl2 + t590_inl2_inl2); */
                    /* c1227 <= (c1223 && c591_inl2_inl2); */
                    /* c1232 <= (c1223 && !c591_inl2_inl2); */
                    /* t594_inl2_inl2 <= (t593_inl2_inl2 << 7); */
                    /* rv_n_inl2_inl24 <= c1227 ? rv_n_inl2_inl23 : (c1223 && !c591_inl2_inl2) ? rv_n_inl2_inl22 : 'bz; */
                    /* t595_inl2_inl2 <= (t592_inl2_inl2 | t594_inl2_inl2); */
                    /* t596_inl2_inl2 <= (rv_n_inl2_inl24 & 127); */
                    /* sub_add_result2_inl22 <= (t595_inl2_inl2 | t596_inl2_inl2); */
                    do_mnist7_mem_state <= do_mnist7_mem_L5_exit104_S0;
                  end else begin
                    /* c1703 <= (c1697 && !c587_inl2_inl2); */
                    /* c1224 <= (c1219 && c643_inl2_inl2); */
                    do_mnist7_mem_state <= do_mnist7_mem_L5_b107_S0;
                  end
                end
              end
            end
          end
        end
      end
      do_mnist7_mem_L5_b91_S0: begin
        i_inl1_inl23 <= 0;
        /* c1222 <= (c1212 && c644_inl1_inl2); */
        /* b_inl1_inl24 <= c1217 ? t569_inl2 : (c1212 && c644_inl1_inl2) ? t570_inl2 : 'bz; */
        /* x_inl1_inl24 <= c1217 ? t570_inl2 : (c1212 && c644_inl1_inl2) ? t569_inl2 : 'bz; */
        /* x_sign_inl1_inl24 <= c1217 ? b_sign_inl24 : (c1212 && c644_inl1_inl2) ? x_sign_inl24 : 'bz; */
        /* rv_n_inl1_inl25 <= (x_inl1_inl24 - b_inl1_inl24); */
        rv_n_inl1_inl26 <= rv_n_inl1_inl25;
        do_mnist7_mem_state <= do_mnist7_mem_L7_fortest92_S0;
      end
      do_mnist7_mem_L5_b107_S0: begin
        i_inl2_inl23 <= 0;
        /* c1228 <= (c1219 && c644_inl2_inl2); */
        /* b_inl2_inl24 <= c1224 ? t577_inl2 : (c1219 && c644_inl2_inl2) ? new_b_n_inl2 : 'bz; */
        /* x_inl2_inl24 <= c1224 ? new_b_n_inl2 : (c1219 && c644_inl2_inl2) ? t577_inl2 : 'bz; */
        /* x_sign_inl2_inl24 <= c1224 ? b_sign_inl24 : (c1219 && c644_inl2_inl2) ? x_sign_inl24 : 'bz; */
        /* rv_n_inl2_inl25 <= (x_inl2_inl24 - b_inl2_inl24); */
        rv_n_inl2_inl26 <= rv_n_inl2_inl25;
        do_mnist7_mem_state <= do_mnist7_mem_L6_fortest108_S0;
      end
      do_mnist7_mem_L5_exit87_S0: begin
        /* c1714 <= (c1695 && !c597_inl1_inl2); */
        /* c1243 <= (c1222 || c1217); */
        /* c1242 <= (c1226 || c1221); */
        /* sub_add_result1_inl25 <= (c1226 || c1221) ? sub_add_result1_inl22 : c1235 ? sub_add_result1_inl23 : (c1222 || c1217) ? 0 : 'bz; */
        do_mnist7_mem_state <= do_mnist7_mem_L5_b89_S0;
      end
      do_mnist7_mem_L5_exit104_S0: begin
        /* c1720 <= (c1703 && !c597_inl2_inl2); */
        /* c1251 <= (c1228 || c1224); */
        /* c1250 <= (c1232 || c1227); */
        /* sub_add_result2_inl25 <= (c1232 || c1227) ? sub_add_result2_inl22 : c1244 ? sub_add_result2_inl23 : (c1228 || c1224) ? 0 : 'bz; */
        do_mnist7_mem_state <= do_mnist7_mem_L5_b89_S0;
      end
      do_mnist7_mem_L5_b89_S0: begin
        /* c1722 <= ((c1694 || c1714) || c1708); */
        /* c1255 <= ((c1242 || c1243) || c1235); */
        /* c1723 <= ((c1702 || c1720) || c1715); */
        /* c1256 <= ((c1250 || c1251) || c1244); */
        /* rv_inl24 <= ((c1242 || c1243) || c1235) ? sub_add_result1_inl25 : ((c1250 || c1251) || c1244) ? sub_add_result2_inl25 : 'bz; */
        /* add_result26 <= rv_inl24; */
        do_mnist7_mem_state <= do_mnist7_mem_L5_exit74_S0;
      end
      do_mnist7_mem_L5_exit74_S0: begin
        _mem_addr <= j6;
        _mem_we <= 1;
        _mem_req <= 1;
        _mem_d <= add_result27;
        /* j7 <= (j6 + 1); */
        /* add_result27 <= c1198 ? t613 : c1202 ? t612 : c1208 ? x_inl24 : c1218 ? x_inl24 : (c1255 || c1256) ? add_result26 : 'bz; */
        j6 <= j7;
        do_mnist7_mem_state <= do_mnist7_mem_L5_exit74_S1;
      end
      do_mnist7_mem_L5_exit74_S1: begin
        _mem_req <= 0;
        do_mnist7_mem_state <= do_mnist7_mem_L5_fortest12_S0;
      end
      do_mnist7_mem_L6_fortest108_S0: begin
        /* c597_inl2_inl2 <= (i_inl2_inl23 < 7); */
        if (c597_inl2_inl2) begin
          /* t598_inl2_inl2 <= (rv_n_inl2_inl26 & 128); */
          /* c1710 <= (c1703 && c597_inl2_inl2); */
          /* c1237 <= ((c1228 || c1224) && c597_inl2_inl2); */
          /* c599_inl2_inl2 <= (t598_inl2_inl2 != 0); */
          if (c599_inl2_inl2) begin
            /* c1715 <= (c1710 && c599_inl2_inl2); */
            /* c1244 <= (c1237 && c599_inl2_inl2); */
            /* t601_inl2_inl2 <= (e_inl2_inl2 - i_inl2_inl23); */
            /* t602_inl2_inl2 <= (t601_inl2_inl2 << 7); */
            /* t600_inl2_inl2 <= x_sign_inl2_inl24 ? 32768 : 0; */
            /* t603_inl2_inl2 <= (t600_inl2_inl2 | t602_inl2_inl2); */
            /* t604_inl2_inl2 <= (rv_n_inl2_inl26 & 127); */
            /* sub_add_result2_inl23 <= (t603_inl2_inl2 | t604_inl2_inl2); */
            do_mnist7_mem_state <= do_mnist7_mem_L5_exit104_S0;
          end else begin
            /* rv_n_inl2_inl27 <= (rv_n_inl2_inl26 << 1); */
            /* i_inl2_inl24 <= (i_inl2_inl23 + 1); */
            i_inl2_inl23 <= i_inl2_inl24;
            rv_n_inl2_inl26 <= rv_n_inl2_inl27;
            /* c1716 <= (c1710 && !c599_inl2_inl2); */
            /* c1245 <= (c1237 && !c599_inl2_inl2); */
            do_mnist7_mem_state <= do_mnist7_mem_L6_fortest108_S0;
          end
        end else begin
          /* c1720 <= (c1703 && !c597_inl2_inl2); */
          /* c1251 <= (c1228 || c1224); */
          /* c1250 <= (c1232 || c1227); */
          /* sub_add_result2_inl25 <= (c1232 || c1227) ? sub_add_result2_inl22 : c1244 ? sub_add_result2_inl23 : (c1228 || c1224) ? 0 : 'bz; */
          do_mnist7_mem_state <= do_mnist7_mem_L5_b89_S0;
        end
      end
      do_mnist7_mem_L7_fortest92_S0: begin
        /* c597_inl1_inl2 <= (i_inl1_inl23 < 7); */
        if (c597_inl1_inl2) begin
          /* t598_inl1_inl2 <= (rv_n_inl1_inl26 & 128); */
          /* c1706 <= (c1695 && c597_inl1_inl2); */
          /* c1231 <= ((c1222 || c1217) && c597_inl1_inl2); */
          /* c599_inl1_inl2 <= (t598_inl1_inl2 != 0); */
          if (c599_inl1_inl2) begin
            /* c1708 <= (c1706 && c599_inl1_inl2); */
            /* c1235 <= (c1231 && c599_inl1_inl2); */
            /* t601_inl1_inl2 <= (e_inl1_inl2 - i_inl1_inl23); */
            /* t602_inl1_inl2 <= (t601_inl1_inl2 << 7); */
            /* t600_inl1_inl2 <= x_sign_inl1_inl24 ? 32768 : 0; */
            /* t603_inl1_inl2 <= (t600_inl1_inl2 | t602_inl1_inl2); */
            /* t604_inl1_inl2 <= (rv_n_inl1_inl26 & 127); */
            /* sub_add_result1_inl23 <= (t603_inl1_inl2 | t604_inl1_inl2); */
            do_mnist7_mem_state <= do_mnist7_mem_L5_exit87_S0;
          end else begin
            /* rv_n_inl1_inl27 <= (rv_n_inl1_inl26 << 1); */
            /* i_inl1_inl24 <= (i_inl1_inl23 + 1); */
            i_inl1_inl23 <= i_inl1_inl24;
            rv_n_inl1_inl26 <= rv_n_inl1_inl27;
            /* c1709 <= (c1706 && !c599_inl1_inl2); */
            /* c1236 <= (c1231 && !c599_inl1_inl2); */
            do_mnist7_mem_state <= do_mnist7_mem_L7_fortest92_S0;
          end
        end else begin
          /* c1714 <= (c1695 && !c597_inl1_inl2); */
          /* c1243 <= (c1222 || c1217); */
          /* c1242 <= (c1226 || c1221); */
          /* sub_add_result1_inl25 <= (c1226 || c1221) ? sub_add_result1_inl22 : c1235 ? sub_add_result1_inl23 : (c1222 || c1217) ? 0 : 'bz; */
          do_mnist7_mem_state <= do_mnist7_mem_L5_b89_S0;
        end
      end
      endcase
    end
  end
  

endmodule

